magic
tech scmos
timestamp 1607511061
<< ab >>
rect -690 70 -668 214
rect -664 70 -534 214
rect -532 144 -500 214
rect -497 144 -467 214
rect -464 144 -407 214
rect -530 141 -498 144
rect -495 141 -407 144
rect -532 70 -500 141
rect -497 70 -467 141
rect -464 70 -407 141
rect -405 70 -383 214
rect -379 70 -249 214
rect -247 144 -215 214
rect -212 144 -182 214
rect -179 144 -122 214
rect -245 140 -213 144
rect -210 140 -122 144
rect -247 139 -213 140
rect -212 139 -122 140
rect -247 70 -215 139
rect -212 70 -182 139
rect -180 70 -122 139
rect -120 70 -98 214
rect -94 70 36 214
rect 38 144 70 214
rect 73 144 103 214
rect 106 144 163 214
rect 40 140 72 144
rect 75 140 163 144
rect 38 139 72 140
rect 73 139 163 140
rect 38 70 70 139
rect 73 70 103 139
rect 105 70 163 139
rect 165 70 187 214
rect 191 70 321 214
rect 323 144 355 214
rect 358 144 388 214
rect 391 144 448 214
rect 325 140 357 144
rect 360 140 448 144
rect 323 139 357 140
rect 358 139 448 140
rect 323 70 355 139
rect 358 70 388 139
rect 390 70 448 139
rect 452 206 508 214
rect 452 170 483 206
rect 484 170 508 206
rect 452 114 508 170
rect 452 70 483 114
rect 484 70 508 114
rect 512 114 568 214
rect 512 78 543 114
rect 544 78 568 114
rect 512 70 568 78
rect 578 70 602 214
rect -690 -280 -668 -136
rect -664 -280 -534 -136
rect -532 -206 -500 -136
rect -497 -206 -467 -136
rect -464 -206 -407 -136
rect -530 -210 -498 -206
rect -495 -210 -407 -206
rect -532 -280 -500 -210
rect -497 -280 -467 -210
rect -464 -280 -407 -210
rect -405 -280 -383 -136
rect -379 -280 -249 -136
rect -247 -206 -215 -136
rect -212 -206 -182 -136
rect -179 -206 -122 -136
rect -245 -210 -213 -206
rect -210 -210 -122 -206
rect -247 -280 -215 -210
rect -212 -280 -182 -210
rect -179 -280 -122 -210
rect -120 -280 -98 -136
rect -94 -280 36 -136
rect 38 -206 70 -136
rect 73 -206 103 -136
rect 106 -206 163 -136
rect 40 -210 72 -206
rect 75 -210 163 -206
rect 38 -280 70 -210
rect 73 -280 103 -210
rect 106 -280 163 -210
rect 165 -280 187 -136
rect 191 -280 321 -136
rect 323 -206 355 -136
rect 358 -206 388 -136
rect 391 -206 448 -136
rect 325 -210 357 -206
rect 360 -210 448 -206
rect 323 -280 355 -210
rect 358 -280 388 -210
rect 391 -280 448 -210
rect 452 -280 540 -136
rect 544 -280 632 -136
<< nwell >>
rect -695 102 607 182
rect -695 -248 637 -168
<< pwell >>
rect -695 182 607 219
rect -695 65 607 102
rect -695 -168 637 -131
rect -695 -285 637 -248
<< poly >>
rect -626 202 -624 207
rect -619 202 -617 207
rect -612 202 -610 207
rect -679 197 -677 202
rect -653 197 -651 202
rect -599 198 -597 203
rect -572 202 -570 207
rect -565 202 -563 207
rect -558 202 -556 207
rect -545 198 -543 203
rect -523 199 -521 203
rect -512 202 -510 207
rect -488 199 -486 203
rect -477 202 -475 207
rect -446 202 -444 207
rect -439 202 -437 207
rect -432 202 -430 207
rect -679 185 -677 188
rect -653 185 -651 188
rect -626 185 -624 189
rect -683 183 -677 185
rect -683 181 -681 183
rect -679 181 -677 183
rect -683 179 -677 181
rect -657 183 -651 185
rect -657 181 -655 183
rect -653 181 -651 183
rect -657 179 -651 181
rect -635 183 -624 185
rect -635 181 -633 183
rect -631 181 -629 183
rect -635 179 -629 181
rect -679 176 -677 179
rect -653 176 -651 179
rect -679 153 -677 158
rect -631 170 -629 179
rect -619 178 -617 189
rect -612 185 -610 189
rect -599 185 -597 189
rect -572 185 -570 189
rect -613 183 -607 185
rect -613 181 -611 183
rect -609 181 -607 183
rect -613 179 -607 181
rect -603 183 -597 185
rect -603 181 -601 183
rect -599 181 -597 183
rect -603 179 -597 181
rect -581 183 -570 185
rect -581 181 -579 183
rect -577 181 -575 183
rect -581 179 -575 181
rect -623 176 -617 178
rect -623 174 -621 176
rect -619 174 -617 176
rect -623 172 -617 174
rect -653 153 -651 158
rect -619 169 -617 172
rect -609 169 -607 179
rect -599 174 -597 179
rect -631 152 -629 157
rect -577 170 -575 179
rect -565 178 -563 189
rect -558 185 -556 189
rect -545 185 -543 189
rect -523 188 -521 191
rect -559 183 -553 185
rect -559 181 -557 183
rect -555 181 -553 183
rect -559 179 -553 181
rect -549 183 -543 185
rect -549 181 -547 183
rect -545 181 -543 183
rect -525 186 -519 188
rect -525 184 -523 186
rect -521 184 -519 186
rect -512 185 -510 194
rect -488 188 -486 191
rect -490 186 -484 188
rect -525 182 -519 184
rect -549 179 -543 181
rect -569 176 -563 178
rect -569 174 -567 176
rect -565 174 -563 176
rect -569 172 -563 174
rect -565 169 -563 172
rect -555 169 -553 179
rect -545 174 -543 179
rect -521 176 -519 182
rect -515 183 -509 185
rect -515 181 -513 183
rect -511 181 -509 183
rect -490 184 -488 186
rect -486 184 -484 186
rect -477 185 -475 194
rect -419 198 -417 203
rect -341 202 -339 207
rect -334 202 -332 207
rect -327 202 -325 207
rect -394 197 -392 202
rect -368 197 -366 202
rect -446 185 -444 189
rect -490 182 -484 184
rect -515 179 -509 181
rect -514 176 -512 179
rect -486 176 -484 182
rect -480 183 -474 185
rect -480 181 -478 183
rect -476 181 -474 183
rect -480 179 -474 181
rect -455 183 -444 185
rect -455 181 -453 183
rect -451 181 -449 183
rect -455 179 -449 181
rect -479 176 -477 179
rect -619 151 -617 156
rect -609 151 -607 156
rect -599 151 -597 156
rect -577 152 -575 157
rect -565 151 -563 156
rect -555 151 -553 156
rect -545 151 -543 156
rect -451 170 -449 179
rect -439 178 -437 189
rect -432 185 -430 189
rect -419 185 -417 189
rect -314 198 -312 203
rect -287 202 -285 207
rect -280 202 -278 207
rect -273 202 -271 207
rect -260 198 -258 203
rect -238 199 -236 203
rect -227 202 -225 207
rect -203 199 -201 203
rect -192 202 -190 207
rect -161 202 -159 207
rect -154 202 -152 207
rect -147 202 -145 207
rect -394 185 -392 188
rect -368 185 -366 188
rect -341 185 -339 189
rect -433 183 -427 185
rect -433 181 -431 183
rect -429 181 -427 183
rect -433 179 -427 181
rect -423 183 -417 185
rect -423 181 -421 183
rect -419 181 -417 183
rect -423 179 -417 181
rect -398 183 -392 185
rect -398 181 -396 183
rect -394 181 -392 183
rect -398 179 -392 181
rect -372 183 -366 185
rect -372 181 -370 183
rect -368 181 -366 183
rect -372 179 -366 181
rect -350 183 -339 185
rect -350 181 -348 183
rect -346 181 -344 183
rect -350 179 -344 181
rect -443 176 -437 178
rect -443 174 -441 176
rect -439 174 -437 176
rect -443 172 -437 174
rect -439 169 -437 172
rect -429 169 -427 179
rect -419 174 -417 179
rect -394 176 -392 179
rect -368 176 -366 179
rect -451 152 -449 157
rect -521 144 -519 148
rect -514 144 -512 148
rect -486 144 -484 148
rect -479 144 -477 148
rect -439 151 -437 156
rect -429 151 -427 156
rect -419 151 -417 156
rect -394 153 -392 158
rect -346 170 -344 179
rect -334 178 -332 189
rect -327 185 -325 189
rect -314 185 -312 189
rect -287 185 -285 189
rect -328 183 -322 185
rect -328 181 -326 183
rect -324 181 -322 183
rect -328 179 -322 181
rect -318 183 -312 185
rect -318 181 -316 183
rect -314 181 -312 183
rect -318 179 -312 181
rect -296 183 -285 185
rect -296 181 -294 183
rect -292 181 -290 183
rect -296 179 -290 181
rect -338 176 -332 178
rect -338 174 -336 176
rect -334 174 -332 176
rect -338 172 -332 174
rect -368 153 -366 158
rect -334 169 -332 172
rect -324 169 -322 179
rect -314 174 -312 179
rect -346 152 -344 157
rect -292 170 -290 179
rect -280 178 -278 189
rect -273 185 -271 189
rect -260 185 -258 189
rect -238 188 -236 191
rect -274 183 -268 185
rect -274 181 -272 183
rect -270 181 -268 183
rect -274 179 -268 181
rect -264 183 -258 185
rect -264 181 -262 183
rect -260 181 -258 183
rect -240 186 -234 188
rect -240 184 -238 186
rect -236 184 -234 186
rect -227 185 -225 194
rect -203 188 -201 191
rect -205 186 -199 188
rect -240 182 -234 184
rect -264 179 -258 181
rect -284 176 -278 178
rect -284 174 -282 176
rect -280 174 -278 176
rect -284 172 -278 174
rect -280 169 -278 172
rect -270 169 -268 179
rect -260 174 -258 179
rect -236 176 -234 182
rect -230 183 -224 185
rect -230 181 -228 183
rect -226 181 -224 183
rect -205 184 -203 186
rect -201 184 -199 186
rect -192 185 -190 194
rect -134 198 -132 203
rect -56 202 -54 207
rect -49 202 -47 207
rect -42 202 -40 207
rect -109 197 -107 202
rect -83 197 -81 202
rect -161 185 -159 189
rect -205 182 -199 184
rect -230 179 -224 181
rect -229 176 -227 179
rect -201 176 -199 182
rect -195 183 -189 185
rect -195 181 -193 183
rect -191 181 -189 183
rect -195 179 -189 181
rect -170 183 -159 185
rect -170 181 -168 183
rect -166 181 -164 183
rect -170 179 -164 181
rect -194 176 -192 179
rect -334 151 -332 156
rect -324 151 -322 156
rect -314 151 -312 156
rect -292 152 -290 157
rect -280 151 -278 156
rect -270 151 -268 156
rect -260 151 -258 156
rect -166 170 -164 179
rect -154 178 -152 189
rect -147 185 -145 189
rect -134 185 -132 189
rect -29 198 -27 203
rect -2 202 0 207
rect 5 202 7 207
rect 12 202 14 207
rect 25 198 27 203
rect 47 199 49 203
rect 58 202 60 207
rect 82 199 84 203
rect 93 202 95 207
rect 124 202 126 207
rect 131 202 133 207
rect 138 202 140 207
rect -109 185 -107 188
rect -83 185 -81 188
rect -56 185 -54 189
rect -148 183 -142 185
rect -148 181 -146 183
rect -144 181 -142 183
rect -148 179 -142 181
rect -138 183 -132 185
rect -138 181 -136 183
rect -134 181 -132 183
rect -138 179 -132 181
rect -113 183 -107 185
rect -113 181 -111 183
rect -109 181 -107 183
rect -113 179 -107 181
rect -87 183 -81 185
rect -87 181 -85 183
rect -83 181 -81 183
rect -87 179 -81 181
rect -65 183 -54 185
rect -65 181 -63 183
rect -61 181 -59 183
rect -65 179 -59 181
rect -158 176 -152 178
rect -158 174 -156 176
rect -154 174 -152 176
rect -158 172 -152 174
rect -154 169 -152 172
rect -144 169 -142 179
rect -134 174 -132 179
rect -109 176 -107 179
rect -83 176 -81 179
rect -166 152 -164 157
rect -236 144 -234 148
rect -229 144 -227 148
rect -201 144 -199 148
rect -194 144 -192 148
rect -154 151 -152 156
rect -144 151 -142 156
rect -134 151 -132 156
rect -109 153 -107 158
rect -61 170 -59 179
rect -49 178 -47 189
rect -42 185 -40 189
rect -29 185 -27 189
rect -2 185 0 189
rect -43 183 -37 185
rect -43 181 -41 183
rect -39 181 -37 183
rect -43 179 -37 181
rect -33 183 -27 185
rect -33 181 -31 183
rect -29 181 -27 183
rect -33 179 -27 181
rect -11 183 0 185
rect -11 181 -9 183
rect -7 181 -5 183
rect -11 179 -5 181
rect -53 176 -47 178
rect -53 174 -51 176
rect -49 174 -47 176
rect -53 172 -47 174
rect -83 153 -81 158
rect -49 169 -47 172
rect -39 169 -37 179
rect -29 174 -27 179
rect -61 152 -59 157
rect -7 170 -5 179
rect 5 178 7 189
rect 12 185 14 189
rect 25 185 27 189
rect 47 188 49 191
rect 11 183 17 185
rect 11 181 13 183
rect 15 181 17 183
rect 11 179 17 181
rect 21 183 27 185
rect 21 181 23 183
rect 25 181 27 183
rect 45 186 51 188
rect 45 184 47 186
rect 49 184 51 186
rect 58 185 60 194
rect 82 188 84 191
rect 80 186 86 188
rect 45 182 51 184
rect 21 179 27 181
rect 1 176 7 178
rect 1 174 3 176
rect 5 174 7 176
rect 1 172 7 174
rect 5 169 7 172
rect 15 169 17 179
rect 25 174 27 179
rect 49 176 51 182
rect 55 183 61 185
rect 55 181 57 183
rect 59 181 61 183
rect 80 184 82 186
rect 84 184 86 186
rect 93 185 95 194
rect 151 198 153 203
rect 229 202 231 207
rect 236 202 238 207
rect 243 202 245 207
rect 176 197 178 202
rect 202 197 204 202
rect 124 185 126 189
rect 80 182 86 184
rect 55 179 61 181
rect 56 176 58 179
rect 84 176 86 182
rect 90 183 96 185
rect 90 181 92 183
rect 94 181 96 183
rect 90 179 96 181
rect 115 183 126 185
rect 115 181 117 183
rect 119 181 121 183
rect 115 179 121 181
rect 91 176 93 179
rect -49 151 -47 156
rect -39 151 -37 156
rect -29 151 -27 156
rect -7 152 -5 157
rect 5 151 7 156
rect 15 151 17 156
rect 25 151 27 156
rect 119 170 121 179
rect 131 178 133 189
rect 138 185 140 189
rect 151 185 153 189
rect 256 198 258 203
rect 283 202 285 207
rect 290 202 292 207
rect 297 202 299 207
rect 310 198 312 203
rect 332 199 334 203
rect 343 202 345 207
rect 367 199 369 203
rect 378 202 380 207
rect 409 202 411 207
rect 416 202 418 207
rect 423 202 425 207
rect 176 185 178 188
rect 202 185 204 188
rect 229 185 231 189
rect 137 183 143 185
rect 137 181 139 183
rect 141 181 143 183
rect 137 179 143 181
rect 147 183 153 185
rect 147 181 149 183
rect 151 181 153 183
rect 147 179 153 181
rect 172 183 178 185
rect 172 181 174 183
rect 176 181 178 183
rect 172 179 178 181
rect 198 183 204 185
rect 198 181 200 183
rect 202 181 204 183
rect 198 179 204 181
rect 220 183 231 185
rect 220 181 222 183
rect 224 181 226 183
rect 220 179 226 181
rect 127 176 133 178
rect 127 174 129 176
rect 131 174 133 176
rect 127 172 133 174
rect 131 169 133 172
rect 141 169 143 179
rect 151 174 153 179
rect 176 176 178 179
rect 202 176 204 179
rect 119 152 121 157
rect 49 144 51 148
rect 56 144 58 148
rect 84 144 86 148
rect 91 144 93 148
rect 131 151 133 156
rect 141 151 143 156
rect 151 151 153 156
rect 176 153 178 158
rect 224 170 226 179
rect 236 178 238 189
rect 243 185 245 189
rect 256 185 258 189
rect 283 185 285 189
rect 242 183 248 185
rect 242 181 244 183
rect 246 181 248 183
rect 242 179 248 181
rect 252 183 258 185
rect 252 181 254 183
rect 256 181 258 183
rect 252 179 258 181
rect 274 183 285 185
rect 274 181 276 183
rect 278 181 280 183
rect 274 179 280 181
rect 232 176 238 178
rect 232 174 234 176
rect 236 174 238 176
rect 232 172 238 174
rect 202 153 204 158
rect 236 169 238 172
rect 246 169 248 179
rect 256 174 258 179
rect 224 152 226 157
rect 278 170 280 179
rect 290 178 292 189
rect 297 185 299 189
rect 310 185 312 189
rect 332 188 334 191
rect 296 183 302 185
rect 296 181 298 183
rect 300 181 302 183
rect 296 179 302 181
rect 306 183 312 185
rect 306 181 308 183
rect 310 181 312 183
rect 330 186 336 188
rect 330 184 332 186
rect 334 184 336 186
rect 343 185 345 194
rect 367 188 369 191
rect 365 186 371 188
rect 330 182 336 184
rect 306 179 312 181
rect 286 176 292 178
rect 286 174 288 176
rect 290 174 292 176
rect 286 172 292 174
rect 290 169 292 172
rect 300 169 302 179
rect 310 174 312 179
rect 334 176 336 182
rect 340 183 346 185
rect 340 181 342 183
rect 344 181 346 183
rect 365 184 367 186
rect 369 184 371 186
rect 378 185 380 194
rect 436 198 438 203
rect 461 198 463 203
rect 474 202 476 207
rect 481 202 483 207
rect 488 202 490 207
rect 521 198 523 203
rect 534 202 536 207
rect 541 202 543 207
rect 548 202 550 207
rect 587 197 589 202
rect 409 185 411 189
rect 365 182 371 184
rect 340 179 346 181
rect 341 176 343 179
rect 369 176 371 182
rect 375 183 381 185
rect 375 181 377 183
rect 379 181 381 183
rect 375 179 381 181
rect 400 183 411 185
rect 400 181 402 183
rect 404 181 406 183
rect 400 179 406 181
rect 376 176 378 179
rect 236 151 238 156
rect 246 151 248 156
rect 256 151 258 156
rect 278 152 280 157
rect 290 151 292 156
rect 300 151 302 156
rect 310 151 312 156
rect 404 170 406 179
rect 416 178 418 189
rect 423 185 425 189
rect 436 185 438 189
rect 422 183 428 185
rect 422 181 424 183
rect 426 181 428 183
rect 422 179 428 181
rect 432 183 438 185
rect 432 181 434 183
rect 436 181 438 183
rect 432 179 438 181
rect 412 176 418 178
rect 412 174 414 176
rect 416 174 418 176
rect 412 172 418 174
rect 416 169 418 172
rect 426 169 428 179
rect 436 174 438 179
rect 461 185 463 189
rect 474 185 476 189
rect 461 183 467 185
rect 461 181 463 183
rect 465 181 467 183
rect 461 179 467 181
rect 471 183 477 185
rect 471 181 473 183
rect 475 181 477 183
rect 471 179 477 181
rect 461 174 463 179
rect 404 152 406 157
rect 471 169 473 179
rect 481 178 483 189
rect 488 185 490 189
rect 521 185 523 189
rect 534 185 536 189
rect 488 183 499 185
rect 493 181 495 183
rect 497 181 499 183
rect 493 179 499 181
rect 521 183 527 185
rect 521 181 523 183
rect 525 181 527 183
rect 521 179 527 181
rect 531 183 537 185
rect 531 181 533 183
rect 535 181 537 183
rect 531 179 537 181
rect 481 176 487 178
rect 481 174 483 176
rect 485 174 487 176
rect 481 172 487 174
rect 481 169 483 172
rect 493 170 495 179
rect 521 174 523 179
rect 334 144 336 148
rect 341 144 343 148
rect 369 144 371 148
rect 376 144 378 148
rect 416 151 418 156
rect 426 151 428 156
rect 436 151 438 156
rect 461 151 463 156
rect 471 151 473 156
rect 481 151 483 156
rect 493 152 495 157
rect 531 169 533 179
rect 541 178 543 189
rect 548 185 550 189
rect 587 185 589 188
rect 548 183 559 185
rect 553 181 555 183
rect 557 181 559 183
rect 553 179 559 181
rect 587 183 593 185
rect 587 181 589 183
rect 591 181 593 183
rect 587 179 593 181
rect 541 176 547 178
rect 541 174 543 176
rect 545 174 547 176
rect 541 172 547 174
rect 541 169 543 172
rect 553 170 555 179
rect 587 176 589 179
rect 521 151 523 156
rect 531 151 533 156
rect 541 151 543 156
rect 553 152 555 157
rect 587 153 589 158
rect -679 126 -677 131
rect -653 126 -651 131
rect -631 127 -629 132
rect -521 136 -519 140
rect -514 136 -512 140
rect -486 136 -484 140
rect -479 136 -477 140
rect -619 128 -617 133
rect -609 128 -607 133
rect -599 128 -597 133
rect -679 105 -677 108
rect -653 105 -651 108
rect -631 105 -629 114
rect -619 112 -617 115
rect -623 110 -617 112
rect -623 108 -621 110
rect -619 108 -617 110
rect -623 106 -617 108
rect -683 103 -677 105
rect -683 101 -681 103
rect -679 101 -677 103
rect -683 99 -677 101
rect -657 103 -651 105
rect -657 101 -655 103
rect -653 101 -651 103
rect -657 99 -651 101
rect -635 103 -629 105
rect -635 101 -633 103
rect -631 101 -629 103
rect -635 99 -624 101
rect -679 96 -677 99
rect -653 96 -651 99
rect -626 95 -624 99
rect -619 95 -617 106
rect -609 105 -607 115
rect -577 127 -575 132
rect -565 128 -563 133
rect -555 128 -553 133
rect -545 128 -543 133
rect -599 105 -597 110
rect -577 105 -575 114
rect -565 112 -563 115
rect -569 110 -563 112
rect -569 108 -567 110
rect -565 108 -563 110
rect -569 106 -563 108
rect -613 103 -607 105
rect -613 101 -611 103
rect -609 101 -607 103
rect -613 99 -607 101
rect -603 103 -597 105
rect -603 101 -601 103
rect -599 101 -597 103
rect -603 99 -597 101
rect -581 103 -575 105
rect -581 101 -579 103
rect -577 101 -575 103
rect -581 99 -570 101
rect -612 95 -610 99
rect -599 95 -597 99
rect -572 95 -570 99
rect -565 95 -563 106
rect -555 105 -553 115
rect -545 105 -543 110
rect -451 127 -449 132
rect -439 128 -437 133
rect -429 128 -427 133
rect -419 128 -417 133
rect -559 103 -553 105
rect -559 101 -557 103
rect -555 101 -553 103
rect -559 99 -553 101
rect -549 103 -543 105
rect -549 101 -547 103
rect -545 101 -543 103
rect -521 102 -519 108
rect -514 105 -512 108
rect -549 99 -543 101
rect -558 95 -556 99
rect -545 95 -543 99
rect -525 100 -519 102
rect -525 98 -523 100
rect -521 98 -519 100
rect -515 103 -509 105
rect -515 101 -513 103
rect -511 101 -509 103
rect -486 102 -484 108
rect -479 105 -477 108
rect -451 105 -449 114
rect -439 112 -437 115
rect -443 110 -437 112
rect -443 108 -441 110
rect -439 108 -437 110
rect -443 106 -437 108
rect -515 99 -509 101
rect -490 100 -484 102
rect -525 96 -519 98
rect -679 82 -677 87
rect -653 82 -651 87
rect -626 77 -624 82
rect -619 77 -617 82
rect -612 77 -610 82
rect -599 81 -597 86
rect -523 93 -521 96
rect -572 77 -570 82
rect -565 77 -563 82
rect -558 77 -556 82
rect -545 81 -543 86
rect -512 90 -510 99
rect -490 98 -488 100
rect -486 98 -484 100
rect -480 103 -474 105
rect -480 101 -478 103
rect -476 101 -474 103
rect -480 99 -474 101
rect -455 103 -449 105
rect -455 101 -453 103
rect -451 101 -449 103
rect -455 99 -444 101
rect -490 96 -484 98
rect -488 93 -486 96
rect -523 81 -521 85
rect -477 90 -475 99
rect -446 95 -444 99
rect -439 95 -437 106
rect -429 105 -427 115
rect -394 126 -392 131
rect -419 105 -417 110
rect -368 126 -366 131
rect -346 127 -344 132
rect -236 136 -234 140
rect -229 136 -227 140
rect -201 136 -199 140
rect -194 136 -192 140
rect -334 128 -332 133
rect -324 128 -322 133
rect -314 128 -312 133
rect -394 105 -392 108
rect -368 105 -366 108
rect -346 105 -344 114
rect -334 112 -332 115
rect -338 110 -332 112
rect -338 108 -336 110
rect -334 108 -332 110
rect -338 106 -332 108
rect -433 103 -427 105
rect -433 101 -431 103
rect -429 101 -427 103
rect -433 99 -427 101
rect -423 103 -417 105
rect -423 101 -421 103
rect -419 101 -417 103
rect -423 99 -417 101
rect -398 103 -392 105
rect -398 101 -396 103
rect -394 101 -392 103
rect -398 99 -392 101
rect -372 103 -366 105
rect -372 101 -370 103
rect -368 101 -366 103
rect -372 99 -366 101
rect -350 103 -344 105
rect -350 101 -348 103
rect -346 101 -344 103
rect -350 99 -339 101
rect -432 95 -430 99
rect -419 95 -417 99
rect -394 96 -392 99
rect -368 96 -366 99
rect -512 77 -510 82
rect -488 81 -486 85
rect -341 95 -339 99
rect -334 95 -332 106
rect -324 105 -322 115
rect -292 127 -290 132
rect -280 128 -278 133
rect -270 128 -268 133
rect -260 128 -258 133
rect -314 105 -312 110
rect -292 105 -290 114
rect -280 112 -278 115
rect -284 110 -278 112
rect -284 108 -282 110
rect -280 108 -278 110
rect -284 106 -278 108
rect -328 103 -322 105
rect -328 101 -326 103
rect -324 101 -322 103
rect -328 99 -322 101
rect -318 103 -312 105
rect -318 101 -316 103
rect -314 101 -312 103
rect -318 99 -312 101
rect -296 103 -290 105
rect -296 101 -294 103
rect -292 101 -290 103
rect -296 99 -285 101
rect -327 95 -325 99
rect -314 95 -312 99
rect -287 95 -285 99
rect -280 95 -278 106
rect -270 105 -268 115
rect -260 105 -258 110
rect -166 127 -164 132
rect -154 128 -152 133
rect -144 128 -142 133
rect -134 128 -132 133
rect -274 103 -268 105
rect -274 101 -272 103
rect -270 101 -268 103
rect -274 99 -268 101
rect -264 103 -258 105
rect -264 101 -262 103
rect -260 101 -258 103
rect -236 102 -234 108
rect -229 105 -227 108
rect -264 99 -258 101
rect -273 95 -271 99
rect -260 95 -258 99
rect -240 100 -234 102
rect -240 98 -238 100
rect -236 98 -234 100
rect -230 103 -224 105
rect -230 101 -228 103
rect -226 101 -224 103
rect -201 102 -199 108
rect -194 105 -192 108
rect -166 105 -164 114
rect -154 112 -152 115
rect -158 110 -152 112
rect -158 108 -156 110
rect -154 108 -152 110
rect -158 106 -152 108
rect -230 99 -224 101
rect -205 100 -199 102
rect -240 96 -234 98
rect -477 77 -475 82
rect -446 77 -444 82
rect -439 77 -437 82
rect -432 77 -430 82
rect -419 81 -417 86
rect -394 82 -392 87
rect -368 82 -366 87
rect -341 77 -339 82
rect -334 77 -332 82
rect -327 77 -325 82
rect -314 81 -312 86
rect -238 93 -236 96
rect -287 77 -285 82
rect -280 77 -278 82
rect -273 77 -271 82
rect -260 81 -258 86
rect -227 90 -225 99
rect -205 98 -203 100
rect -201 98 -199 100
rect -195 103 -189 105
rect -195 101 -193 103
rect -191 101 -189 103
rect -195 99 -189 101
rect -170 103 -164 105
rect -170 101 -168 103
rect -166 101 -164 103
rect -170 99 -159 101
rect -205 96 -199 98
rect -203 93 -201 96
rect -238 81 -236 85
rect -192 90 -190 99
rect -161 95 -159 99
rect -154 95 -152 106
rect -144 105 -142 115
rect -109 126 -107 131
rect -134 105 -132 110
rect -83 126 -81 131
rect -61 127 -59 132
rect 49 136 51 140
rect 56 136 58 140
rect 84 136 86 140
rect 91 136 93 140
rect -49 128 -47 133
rect -39 128 -37 133
rect -29 128 -27 133
rect -109 105 -107 108
rect -83 105 -81 108
rect -61 105 -59 114
rect -49 112 -47 115
rect -53 110 -47 112
rect -53 108 -51 110
rect -49 108 -47 110
rect -53 106 -47 108
rect -148 103 -142 105
rect -148 101 -146 103
rect -144 101 -142 103
rect -148 99 -142 101
rect -138 103 -132 105
rect -138 101 -136 103
rect -134 101 -132 103
rect -138 99 -132 101
rect -113 103 -107 105
rect -113 101 -111 103
rect -109 101 -107 103
rect -113 99 -107 101
rect -87 103 -81 105
rect -87 101 -85 103
rect -83 101 -81 103
rect -87 99 -81 101
rect -65 103 -59 105
rect -65 101 -63 103
rect -61 101 -59 103
rect -65 99 -54 101
rect -147 95 -145 99
rect -134 95 -132 99
rect -109 96 -107 99
rect -83 96 -81 99
rect -227 77 -225 82
rect -203 81 -201 85
rect -56 95 -54 99
rect -49 95 -47 106
rect -39 105 -37 115
rect -7 127 -5 132
rect 5 128 7 133
rect 15 128 17 133
rect 25 128 27 133
rect -29 105 -27 110
rect -7 105 -5 114
rect 5 112 7 115
rect 1 110 7 112
rect 1 108 3 110
rect 5 108 7 110
rect 1 106 7 108
rect -43 103 -37 105
rect -43 101 -41 103
rect -39 101 -37 103
rect -43 99 -37 101
rect -33 103 -27 105
rect -33 101 -31 103
rect -29 101 -27 103
rect -33 99 -27 101
rect -11 103 -5 105
rect -11 101 -9 103
rect -7 101 -5 103
rect -11 99 0 101
rect -42 95 -40 99
rect -29 95 -27 99
rect -2 95 0 99
rect 5 95 7 106
rect 15 105 17 115
rect 25 105 27 110
rect 119 127 121 132
rect 131 128 133 133
rect 141 128 143 133
rect 151 128 153 133
rect 11 103 17 105
rect 11 101 13 103
rect 15 101 17 103
rect 11 99 17 101
rect 21 103 27 105
rect 21 101 23 103
rect 25 101 27 103
rect 49 102 51 108
rect 56 105 58 108
rect 21 99 27 101
rect 12 95 14 99
rect 25 95 27 99
rect 45 100 51 102
rect 45 98 47 100
rect 49 98 51 100
rect 55 103 61 105
rect 55 101 57 103
rect 59 101 61 103
rect 84 102 86 108
rect 91 105 93 108
rect 119 105 121 114
rect 131 112 133 115
rect 127 110 133 112
rect 127 108 129 110
rect 131 108 133 110
rect 127 106 133 108
rect 55 99 61 101
rect 80 100 86 102
rect 45 96 51 98
rect -192 77 -190 82
rect -161 77 -159 82
rect -154 77 -152 82
rect -147 77 -145 82
rect -134 81 -132 86
rect -109 82 -107 87
rect -83 82 -81 87
rect -56 77 -54 82
rect -49 77 -47 82
rect -42 77 -40 82
rect -29 81 -27 86
rect 47 93 49 96
rect -2 77 0 82
rect 5 77 7 82
rect 12 77 14 82
rect 25 81 27 86
rect 58 90 60 99
rect 80 98 82 100
rect 84 98 86 100
rect 90 103 96 105
rect 90 101 92 103
rect 94 101 96 103
rect 90 99 96 101
rect 115 103 121 105
rect 115 101 117 103
rect 119 101 121 103
rect 115 99 126 101
rect 80 96 86 98
rect 82 93 84 96
rect 47 81 49 85
rect 93 90 95 99
rect 124 95 126 99
rect 131 95 133 106
rect 141 105 143 115
rect 176 126 178 131
rect 151 105 153 110
rect 202 126 204 131
rect 224 127 226 132
rect 334 136 336 140
rect 341 136 343 140
rect 369 136 371 140
rect 376 136 378 140
rect 236 128 238 133
rect 246 128 248 133
rect 256 128 258 133
rect 176 105 178 108
rect 202 105 204 108
rect 224 105 226 114
rect 236 112 238 115
rect 232 110 238 112
rect 232 108 234 110
rect 236 108 238 110
rect 232 106 238 108
rect 137 103 143 105
rect 137 101 139 103
rect 141 101 143 103
rect 137 99 143 101
rect 147 103 153 105
rect 147 101 149 103
rect 151 101 153 103
rect 147 99 153 101
rect 172 103 178 105
rect 172 101 174 103
rect 176 101 178 103
rect 172 99 178 101
rect 198 103 204 105
rect 198 101 200 103
rect 202 101 204 103
rect 198 99 204 101
rect 220 103 226 105
rect 220 101 222 103
rect 224 101 226 103
rect 220 99 231 101
rect 138 95 140 99
rect 151 95 153 99
rect 176 96 178 99
rect 202 96 204 99
rect 58 77 60 82
rect 82 81 84 85
rect 229 95 231 99
rect 236 95 238 106
rect 246 105 248 115
rect 278 127 280 132
rect 290 128 292 133
rect 300 128 302 133
rect 310 128 312 133
rect 256 105 258 110
rect 278 105 280 114
rect 290 112 292 115
rect 286 110 292 112
rect 286 108 288 110
rect 290 108 292 110
rect 286 106 292 108
rect 242 103 248 105
rect 242 101 244 103
rect 246 101 248 103
rect 242 99 248 101
rect 252 103 258 105
rect 252 101 254 103
rect 256 101 258 103
rect 252 99 258 101
rect 274 103 280 105
rect 274 101 276 103
rect 278 101 280 103
rect 274 99 285 101
rect 243 95 245 99
rect 256 95 258 99
rect 283 95 285 99
rect 290 95 292 106
rect 300 105 302 115
rect 310 105 312 110
rect 404 127 406 132
rect 416 128 418 133
rect 426 128 428 133
rect 436 128 438 133
rect 461 128 463 133
rect 471 128 473 133
rect 481 128 483 133
rect 296 103 302 105
rect 296 101 298 103
rect 300 101 302 103
rect 296 99 302 101
rect 306 103 312 105
rect 306 101 308 103
rect 310 101 312 103
rect 334 102 336 108
rect 341 105 343 108
rect 306 99 312 101
rect 297 95 299 99
rect 310 95 312 99
rect 330 100 336 102
rect 330 98 332 100
rect 334 98 336 100
rect 340 103 346 105
rect 340 101 342 103
rect 344 101 346 103
rect 369 102 371 108
rect 376 105 378 108
rect 404 105 406 114
rect 416 112 418 115
rect 412 110 418 112
rect 412 108 414 110
rect 416 108 418 110
rect 412 106 418 108
rect 340 99 346 101
rect 365 100 371 102
rect 330 96 336 98
rect 93 77 95 82
rect 124 77 126 82
rect 131 77 133 82
rect 138 77 140 82
rect 151 81 153 86
rect 176 82 178 87
rect 202 82 204 87
rect 229 77 231 82
rect 236 77 238 82
rect 243 77 245 82
rect 256 81 258 86
rect 332 93 334 96
rect 283 77 285 82
rect 290 77 292 82
rect 297 77 299 82
rect 310 81 312 86
rect 343 90 345 99
rect 365 98 367 100
rect 369 98 371 100
rect 375 103 381 105
rect 375 101 377 103
rect 379 101 381 103
rect 375 99 381 101
rect 400 103 406 105
rect 400 101 402 103
rect 404 101 406 103
rect 400 99 411 101
rect 365 96 371 98
rect 367 93 369 96
rect 332 81 334 85
rect 378 90 380 99
rect 409 95 411 99
rect 416 95 418 106
rect 426 105 428 115
rect 493 127 495 132
rect 521 128 523 133
rect 531 128 533 133
rect 541 128 543 133
rect 436 105 438 110
rect 422 103 428 105
rect 422 101 424 103
rect 426 101 428 103
rect 422 99 428 101
rect 432 103 438 105
rect 432 101 434 103
rect 436 101 438 103
rect 432 99 438 101
rect 423 95 425 99
rect 436 95 438 99
rect 461 105 463 110
rect 471 105 473 115
rect 481 112 483 115
rect 481 110 487 112
rect 481 108 483 110
rect 485 108 487 110
rect 481 106 487 108
rect 461 103 467 105
rect 461 101 463 103
rect 465 101 467 103
rect 461 99 467 101
rect 471 103 477 105
rect 471 101 473 103
rect 475 101 477 103
rect 471 99 477 101
rect 461 95 463 99
rect 474 95 476 99
rect 481 95 483 106
rect 493 105 495 114
rect 553 127 555 132
rect 521 105 523 110
rect 531 105 533 115
rect 541 112 543 115
rect 587 126 589 131
rect 541 110 547 112
rect 541 108 543 110
rect 545 108 547 110
rect 541 106 547 108
rect 493 103 499 105
rect 493 101 495 103
rect 497 101 499 103
rect 488 99 499 101
rect 521 103 527 105
rect 521 101 523 103
rect 525 101 527 103
rect 521 99 527 101
rect 531 103 537 105
rect 531 101 533 103
rect 535 101 537 103
rect 531 99 537 101
rect 488 95 490 99
rect 521 95 523 99
rect 534 95 536 99
rect 541 95 543 106
rect 553 105 555 114
rect 587 105 589 108
rect 553 103 559 105
rect 553 101 555 103
rect 557 101 559 103
rect 548 99 559 101
rect 587 103 593 105
rect 587 101 589 103
rect 591 101 593 103
rect 587 99 593 101
rect 548 95 550 99
rect 587 96 589 99
rect 343 77 345 82
rect 367 81 369 85
rect 378 77 380 82
rect 409 77 411 82
rect 416 77 418 82
rect 423 77 425 82
rect 436 81 438 86
rect 461 81 463 86
rect 474 77 476 82
rect 481 77 483 82
rect 488 77 490 82
rect 521 81 523 86
rect 587 82 589 87
rect 534 77 536 82
rect 541 77 543 82
rect 548 77 550 82
rect -626 -148 -624 -143
rect -619 -148 -617 -143
rect -612 -148 -610 -143
rect -679 -153 -677 -148
rect -653 -153 -651 -148
rect -599 -152 -597 -147
rect -572 -148 -570 -143
rect -565 -148 -563 -143
rect -558 -148 -556 -143
rect -545 -152 -543 -147
rect -523 -151 -521 -147
rect -512 -148 -510 -143
rect -488 -151 -486 -147
rect -477 -148 -475 -143
rect -446 -148 -444 -143
rect -439 -148 -437 -143
rect -432 -148 -430 -143
rect -679 -165 -677 -162
rect -653 -165 -651 -162
rect -626 -165 -624 -161
rect -683 -167 -677 -165
rect -683 -169 -681 -167
rect -679 -169 -677 -167
rect -683 -171 -677 -169
rect -657 -167 -651 -165
rect -657 -169 -655 -167
rect -653 -169 -651 -167
rect -657 -171 -651 -169
rect -635 -167 -624 -165
rect -635 -169 -633 -167
rect -631 -169 -629 -167
rect -635 -171 -629 -169
rect -679 -174 -677 -171
rect -653 -174 -651 -171
rect -679 -197 -677 -192
rect -631 -180 -629 -171
rect -619 -172 -617 -161
rect -612 -165 -610 -161
rect -599 -165 -597 -161
rect -572 -165 -570 -161
rect -613 -167 -607 -165
rect -613 -169 -611 -167
rect -609 -169 -607 -167
rect -613 -171 -607 -169
rect -603 -167 -597 -165
rect -603 -169 -601 -167
rect -599 -169 -597 -167
rect -603 -171 -597 -169
rect -581 -167 -570 -165
rect -581 -169 -579 -167
rect -577 -169 -575 -167
rect -581 -171 -575 -169
rect -623 -174 -617 -172
rect -623 -176 -621 -174
rect -619 -176 -617 -174
rect -623 -178 -617 -176
rect -653 -197 -651 -192
rect -619 -181 -617 -178
rect -609 -181 -607 -171
rect -599 -176 -597 -171
rect -631 -198 -629 -193
rect -577 -180 -575 -171
rect -565 -172 -563 -161
rect -558 -165 -556 -161
rect -545 -165 -543 -161
rect -523 -162 -521 -159
rect -559 -167 -553 -165
rect -559 -169 -557 -167
rect -555 -169 -553 -167
rect -559 -171 -553 -169
rect -549 -167 -543 -165
rect -549 -169 -547 -167
rect -545 -169 -543 -167
rect -525 -164 -519 -162
rect -525 -166 -523 -164
rect -521 -166 -519 -164
rect -512 -165 -510 -156
rect -488 -162 -486 -159
rect -490 -164 -484 -162
rect -525 -168 -519 -166
rect -549 -171 -543 -169
rect -569 -174 -563 -172
rect -569 -176 -567 -174
rect -565 -176 -563 -174
rect -569 -178 -563 -176
rect -565 -181 -563 -178
rect -555 -181 -553 -171
rect -545 -176 -543 -171
rect -521 -174 -519 -168
rect -515 -167 -509 -165
rect -515 -169 -513 -167
rect -511 -169 -509 -167
rect -490 -166 -488 -164
rect -486 -166 -484 -164
rect -477 -165 -475 -156
rect -419 -152 -417 -147
rect -341 -148 -339 -143
rect -334 -148 -332 -143
rect -327 -148 -325 -143
rect -394 -153 -392 -148
rect -368 -153 -366 -148
rect -446 -165 -444 -161
rect -490 -168 -484 -166
rect -515 -171 -509 -169
rect -514 -174 -512 -171
rect -486 -174 -484 -168
rect -480 -167 -474 -165
rect -480 -169 -478 -167
rect -476 -169 -474 -167
rect -480 -171 -474 -169
rect -455 -167 -444 -165
rect -455 -169 -453 -167
rect -451 -169 -449 -167
rect -455 -171 -449 -169
rect -479 -174 -477 -171
rect -619 -199 -617 -194
rect -609 -199 -607 -194
rect -599 -199 -597 -194
rect -577 -198 -575 -193
rect -565 -199 -563 -194
rect -555 -199 -553 -194
rect -545 -199 -543 -194
rect -451 -180 -449 -171
rect -439 -172 -437 -161
rect -432 -165 -430 -161
rect -419 -165 -417 -161
rect -314 -152 -312 -147
rect -287 -148 -285 -143
rect -280 -148 -278 -143
rect -273 -148 -271 -143
rect -260 -152 -258 -147
rect -238 -151 -236 -147
rect -227 -148 -225 -143
rect -203 -151 -201 -147
rect -192 -148 -190 -143
rect -161 -148 -159 -143
rect -154 -148 -152 -143
rect -147 -148 -145 -143
rect -394 -165 -392 -162
rect -368 -165 -366 -162
rect -341 -165 -339 -161
rect -433 -167 -427 -165
rect -433 -169 -431 -167
rect -429 -169 -427 -167
rect -433 -171 -427 -169
rect -423 -167 -417 -165
rect -423 -169 -421 -167
rect -419 -169 -417 -167
rect -423 -171 -417 -169
rect -398 -167 -392 -165
rect -398 -169 -396 -167
rect -394 -169 -392 -167
rect -398 -171 -392 -169
rect -372 -167 -366 -165
rect -372 -169 -370 -167
rect -368 -169 -366 -167
rect -372 -171 -366 -169
rect -350 -167 -339 -165
rect -350 -169 -348 -167
rect -346 -169 -344 -167
rect -350 -171 -344 -169
rect -443 -174 -437 -172
rect -443 -176 -441 -174
rect -439 -176 -437 -174
rect -443 -178 -437 -176
rect -439 -181 -437 -178
rect -429 -181 -427 -171
rect -419 -176 -417 -171
rect -394 -174 -392 -171
rect -368 -174 -366 -171
rect -451 -198 -449 -193
rect -521 -206 -519 -202
rect -514 -206 -512 -202
rect -486 -206 -484 -202
rect -479 -206 -477 -202
rect -439 -199 -437 -194
rect -429 -199 -427 -194
rect -419 -199 -417 -194
rect -394 -197 -392 -192
rect -346 -180 -344 -171
rect -334 -172 -332 -161
rect -327 -165 -325 -161
rect -314 -165 -312 -161
rect -287 -165 -285 -161
rect -328 -167 -322 -165
rect -328 -169 -326 -167
rect -324 -169 -322 -167
rect -328 -171 -322 -169
rect -318 -167 -312 -165
rect -318 -169 -316 -167
rect -314 -169 -312 -167
rect -318 -171 -312 -169
rect -296 -167 -285 -165
rect -296 -169 -294 -167
rect -292 -169 -290 -167
rect -296 -171 -290 -169
rect -338 -174 -332 -172
rect -338 -176 -336 -174
rect -334 -176 -332 -174
rect -338 -178 -332 -176
rect -368 -197 -366 -192
rect -334 -181 -332 -178
rect -324 -181 -322 -171
rect -314 -176 -312 -171
rect -346 -198 -344 -193
rect -292 -180 -290 -171
rect -280 -172 -278 -161
rect -273 -165 -271 -161
rect -260 -165 -258 -161
rect -238 -162 -236 -159
rect -274 -167 -268 -165
rect -274 -169 -272 -167
rect -270 -169 -268 -167
rect -274 -171 -268 -169
rect -264 -167 -258 -165
rect -264 -169 -262 -167
rect -260 -169 -258 -167
rect -240 -164 -234 -162
rect -240 -166 -238 -164
rect -236 -166 -234 -164
rect -227 -165 -225 -156
rect -203 -162 -201 -159
rect -205 -164 -199 -162
rect -240 -168 -234 -166
rect -264 -171 -258 -169
rect -284 -174 -278 -172
rect -284 -176 -282 -174
rect -280 -176 -278 -174
rect -284 -178 -278 -176
rect -280 -181 -278 -178
rect -270 -181 -268 -171
rect -260 -176 -258 -171
rect -236 -174 -234 -168
rect -230 -167 -224 -165
rect -230 -169 -228 -167
rect -226 -169 -224 -167
rect -205 -166 -203 -164
rect -201 -166 -199 -164
rect -192 -165 -190 -156
rect -134 -152 -132 -147
rect -56 -148 -54 -143
rect -49 -148 -47 -143
rect -42 -148 -40 -143
rect -109 -153 -107 -148
rect -83 -153 -81 -148
rect -161 -165 -159 -161
rect -205 -168 -199 -166
rect -230 -171 -224 -169
rect -229 -174 -227 -171
rect -201 -174 -199 -168
rect -195 -167 -189 -165
rect -195 -169 -193 -167
rect -191 -169 -189 -167
rect -195 -171 -189 -169
rect -170 -167 -159 -165
rect -170 -169 -168 -167
rect -166 -169 -164 -167
rect -170 -171 -164 -169
rect -194 -174 -192 -171
rect -334 -199 -332 -194
rect -324 -199 -322 -194
rect -314 -199 -312 -194
rect -292 -198 -290 -193
rect -280 -199 -278 -194
rect -270 -199 -268 -194
rect -260 -199 -258 -194
rect -166 -180 -164 -171
rect -154 -172 -152 -161
rect -147 -165 -145 -161
rect -134 -165 -132 -161
rect -29 -152 -27 -147
rect -2 -148 0 -143
rect 5 -148 7 -143
rect 12 -148 14 -143
rect 25 -152 27 -147
rect 47 -151 49 -147
rect 58 -148 60 -143
rect 82 -151 84 -147
rect 93 -148 95 -143
rect 124 -148 126 -143
rect 131 -148 133 -143
rect 138 -148 140 -143
rect -109 -165 -107 -162
rect -83 -165 -81 -162
rect -56 -165 -54 -161
rect -148 -167 -142 -165
rect -148 -169 -146 -167
rect -144 -169 -142 -167
rect -148 -171 -142 -169
rect -138 -167 -132 -165
rect -138 -169 -136 -167
rect -134 -169 -132 -167
rect -138 -171 -132 -169
rect -113 -167 -107 -165
rect -113 -169 -111 -167
rect -109 -169 -107 -167
rect -113 -171 -107 -169
rect -87 -167 -81 -165
rect -87 -169 -85 -167
rect -83 -169 -81 -167
rect -87 -171 -81 -169
rect -65 -167 -54 -165
rect -65 -169 -63 -167
rect -61 -169 -59 -167
rect -65 -171 -59 -169
rect -158 -174 -152 -172
rect -158 -176 -156 -174
rect -154 -176 -152 -174
rect -158 -178 -152 -176
rect -154 -181 -152 -178
rect -144 -181 -142 -171
rect -134 -176 -132 -171
rect -109 -174 -107 -171
rect -83 -174 -81 -171
rect -166 -198 -164 -193
rect -236 -206 -234 -202
rect -229 -206 -227 -202
rect -201 -206 -199 -202
rect -194 -206 -192 -202
rect -154 -199 -152 -194
rect -144 -199 -142 -194
rect -134 -199 -132 -194
rect -109 -197 -107 -192
rect -61 -180 -59 -171
rect -49 -172 -47 -161
rect -42 -165 -40 -161
rect -29 -165 -27 -161
rect -2 -165 0 -161
rect -43 -167 -37 -165
rect -43 -169 -41 -167
rect -39 -169 -37 -167
rect -43 -171 -37 -169
rect -33 -167 -27 -165
rect -33 -169 -31 -167
rect -29 -169 -27 -167
rect -33 -171 -27 -169
rect -11 -167 0 -165
rect -11 -169 -9 -167
rect -7 -169 -5 -167
rect -11 -171 -5 -169
rect -53 -174 -47 -172
rect -53 -176 -51 -174
rect -49 -176 -47 -174
rect -53 -178 -47 -176
rect -83 -197 -81 -192
rect -49 -181 -47 -178
rect -39 -181 -37 -171
rect -29 -176 -27 -171
rect -61 -198 -59 -193
rect -7 -180 -5 -171
rect 5 -172 7 -161
rect 12 -165 14 -161
rect 25 -165 27 -161
rect 47 -162 49 -159
rect 11 -167 17 -165
rect 11 -169 13 -167
rect 15 -169 17 -167
rect 11 -171 17 -169
rect 21 -167 27 -165
rect 21 -169 23 -167
rect 25 -169 27 -167
rect 45 -164 51 -162
rect 45 -166 47 -164
rect 49 -166 51 -164
rect 58 -165 60 -156
rect 82 -162 84 -159
rect 80 -164 86 -162
rect 45 -168 51 -166
rect 21 -171 27 -169
rect 1 -174 7 -172
rect 1 -176 3 -174
rect 5 -176 7 -174
rect 1 -178 7 -176
rect 5 -181 7 -178
rect 15 -181 17 -171
rect 25 -176 27 -171
rect 49 -174 51 -168
rect 55 -167 61 -165
rect 55 -169 57 -167
rect 59 -169 61 -167
rect 80 -166 82 -164
rect 84 -166 86 -164
rect 93 -165 95 -156
rect 151 -152 153 -147
rect 229 -148 231 -143
rect 236 -148 238 -143
rect 243 -148 245 -143
rect 176 -153 178 -148
rect 202 -153 204 -148
rect 124 -165 126 -161
rect 80 -168 86 -166
rect 55 -171 61 -169
rect 56 -174 58 -171
rect 84 -174 86 -168
rect 90 -167 96 -165
rect 90 -169 92 -167
rect 94 -169 96 -167
rect 90 -171 96 -169
rect 115 -167 126 -165
rect 115 -169 117 -167
rect 119 -169 121 -167
rect 115 -171 121 -169
rect 91 -174 93 -171
rect -49 -199 -47 -194
rect -39 -199 -37 -194
rect -29 -199 -27 -194
rect -7 -198 -5 -193
rect 5 -199 7 -194
rect 15 -199 17 -194
rect 25 -199 27 -194
rect 119 -180 121 -171
rect 131 -172 133 -161
rect 138 -165 140 -161
rect 151 -165 153 -161
rect 256 -152 258 -147
rect 283 -148 285 -143
rect 290 -148 292 -143
rect 297 -148 299 -143
rect 310 -152 312 -147
rect 332 -151 334 -147
rect 343 -148 345 -143
rect 367 -151 369 -147
rect 378 -148 380 -143
rect 409 -148 411 -143
rect 416 -148 418 -143
rect 423 -148 425 -143
rect 176 -165 178 -162
rect 202 -165 204 -162
rect 229 -165 231 -161
rect 137 -167 143 -165
rect 137 -169 139 -167
rect 141 -169 143 -167
rect 137 -171 143 -169
rect 147 -167 153 -165
rect 147 -169 149 -167
rect 151 -169 153 -167
rect 147 -171 153 -169
rect 172 -167 178 -165
rect 172 -169 174 -167
rect 176 -169 178 -167
rect 172 -171 178 -169
rect 198 -167 204 -165
rect 198 -169 200 -167
rect 202 -169 204 -167
rect 198 -171 204 -169
rect 220 -167 231 -165
rect 220 -169 222 -167
rect 224 -169 226 -167
rect 220 -171 226 -169
rect 127 -174 133 -172
rect 127 -176 129 -174
rect 131 -176 133 -174
rect 127 -178 133 -176
rect 131 -181 133 -178
rect 141 -181 143 -171
rect 151 -176 153 -171
rect 176 -174 178 -171
rect 202 -174 204 -171
rect 119 -198 121 -193
rect 49 -206 51 -202
rect 56 -206 58 -202
rect 84 -206 86 -202
rect 91 -206 93 -202
rect 131 -199 133 -194
rect 141 -199 143 -194
rect 151 -199 153 -194
rect 176 -197 178 -192
rect 224 -180 226 -171
rect 236 -172 238 -161
rect 243 -165 245 -161
rect 256 -165 258 -161
rect 283 -165 285 -161
rect 242 -167 248 -165
rect 242 -169 244 -167
rect 246 -169 248 -167
rect 242 -171 248 -169
rect 252 -167 258 -165
rect 252 -169 254 -167
rect 256 -169 258 -167
rect 252 -171 258 -169
rect 274 -167 285 -165
rect 274 -169 276 -167
rect 278 -169 280 -167
rect 274 -171 280 -169
rect 232 -174 238 -172
rect 232 -176 234 -174
rect 236 -176 238 -174
rect 232 -178 238 -176
rect 202 -197 204 -192
rect 236 -181 238 -178
rect 246 -181 248 -171
rect 256 -176 258 -171
rect 224 -198 226 -193
rect 278 -180 280 -171
rect 290 -172 292 -161
rect 297 -165 299 -161
rect 310 -165 312 -161
rect 332 -162 334 -159
rect 296 -167 302 -165
rect 296 -169 298 -167
rect 300 -169 302 -167
rect 296 -171 302 -169
rect 306 -167 312 -165
rect 306 -169 308 -167
rect 310 -169 312 -167
rect 330 -164 336 -162
rect 330 -166 332 -164
rect 334 -166 336 -164
rect 343 -165 345 -156
rect 367 -162 369 -159
rect 365 -164 371 -162
rect 330 -168 336 -166
rect 306 -171 312 -169
rect 286 -174 292 -172
rect 286 -176 288 -174
rect 290 -176 292 -174
rect 286 -178 292 -176
rect 290 -181 292 -178
rect 300 -181 302 -171
rect 310 -176 312 -171
rect 334 -174 336 -168
rect 340 -167 346 -165
rect 340 -169 342 -167
rect 344 -169 346 -167
rect 365 -166 367 -164
rect 369 -166 371 -164
rect 378 -165 380 -156
rect 436 -152 438 -147
rect 485 -148 487 -143
rect 495 -148 497 -143
rect 507 -148 509 -143
rect 517 -148 519 -143
rect 529 -148 531 -143
rect 475 -159 481 -157
rect 475 -161 477 -159
rect 479 -161 481 -159
rect 409 -165 411 -161
rect 365 -168 371 -166
rect 340 -171 346 -169
rect 341 -174 343 -171
rect 369 -174 371 -168
rect 375 -167 381 -165
rect 375 -169 377 -167
rect 379 -169 381 -167
rect 375 -171 381 -169
rect 400 -167 411 -165
rect 400 -169 402 -167
rect 404 -169 406 -167
rect 400 -171 406 -169
rect 376 -174 378 -171
rect 236 -199 238 -194
rect 246 -199 248 -194
rect 256 -199 258 -194
rect 278 -198 280 -193
rect 290 -199 292 -194
rect 300 -199 302 -194
rect 310 -199 312 -194
rect 404 -180 406 -171
rect 416 -172 418 -161
rect 423 -165 425 -161
rect 436 -165 438 -161
rect 475 -163 481 -161
rect 422 -167 428 -165
rect 422 -169 424 -167
rect 426 -169 428 -167
rect 422 -171 428 -169
rect 432 -167 438 -165
rect 432 -169 434 -167
rect 436 -169 438 -167
rect 432 -171 438 -169
rect 412 -174 418 -172
rect 412 -176 414 -174
rect 416 -176 418 -174
rect 412 -178 418 -176
rect 416 -181 418 -178
rect 426 -181 428 -171
rect 436 -176 438 -171
rect 469 -169 475 -167
rect 469 -171 471 -169
rect 473 -171 475 -169
rect 469 -173 475 -171
rect 459 -175 465 -173
rect 404 -198 406 -193
rect 459 -177 461 -175
rect 463 -177 465 -175
rect 459 -179 467 -177
rect 465 -182 467 -179
rect 472 -182 474 -173
rect 479 -182 481 -163
rect 485 -173 487 -154
rect 495 -157 497 -154
rect 491 -159 497 -157
rect 491 -161 493 -159
rect 495 -161 497 -159
rect 507 -161 509 -154
rect 491 -163 497 -161
rect 495 -171 497 -163
rect 501 -163 509 -161
rect 501 -165 503 -163
rect 505 -165 509 -163
rect 501 -167 512 -165
rect 495 -173 505 -171
rect 485 -175 491 -173
rect 485 -177 487 -175
rect 489 -177 491 -175
rect 485 -179 498 -177
rect 486 -182 488 -179
rect 496 -182 498 -179
rect 503 -182 505 -173
rect 510 -182 512 -167
rect 517 -171 519 -154
rect 529 -160 531 -157
rect 577 -148 579 -143
rect 587 -148 589 -143
rect 599 -148 601 -143
rect 609 -148 611 -143
rect 621 -148 623 -143
rect 567 -159 573 -157
rect 525 -162 531 -160
rect 525 -164 527 -162
rect 529 -164 531 -162
rect 567 -161 569 -159
rect 571 -161 573 -159
rect 567 -163 573 -161
rect 525 -166 531 -164
rect 516 -173 522 -171
rect 516 -175 518 -173
rect 520 -175 522 -173
rect 529 -174 531 -166
rect 561 -169 567 -167
rect 561 -171 563 -169
rect 565 -171 567 -169
rect 561 -173 567 -171
rect 516 -177 522 -175
rect 517 -182 519 -177
rect 334 -206 336 -202
rect 341 -206 343 -202
rect 369 -206 371 -202
rect 376 -206 378 -202
rect 416 -199 418 -194
rect 426 -199 428 -194
rect 436 -199 438 -194
rect 551 -175 557 -173
rect 551 -177 553 -175
rect 555 -177 557 -175
rect 551 -179 559 -177
rect 557 -182 559 -179
rect 564 -182 566 -173
rect 571 -182 573 -163
rect 577 -173 579 -154
rect 587 -157 589 -154
rect 583 -159 589 -157
rect 583 -161 585 -159
rect 587 -161 589 -159
rect 599 -161 601 -154
rect 583 -163 589 -161
rect 587 -171 589 -163
rect 593 -163 601 -161
rect 593 -165 595 -163
rect 597 -165 601 -163
rect 593 -167 604 -165
rect 587 -173 597 -171
rect 577 -175 583 -173
rect 577 -177 579 -175
rect 581 -177 583 -175
rect 577 -179 590 -177
rect 578 -182 580 -179
rect 588 -182 590 -179
rect 595 -182 597 -173
rect 602 -182 604 -167
rect 609 -171 611 -154
rect 621 -160 623 -157
rect 617 -162 623 -160
rect 617 -164 619 -162
rect 621 -164 623 -162
rect 617 -166 623 -164
rect 608 -173 614 -171
rect 608 -175 610 -173
rect 612 -175 614 -173
rect 621 -174 623 -166
rect 608 -177 614 -175
rect 609 -182 611 -177
rect 529 -197 531 -192
rect 465 -205 467 -200
rect 472 -205 474 -200
rect 479 -205 481 -200
rect 486 -205 488 -200
rect 496 -205 498 -200
rect 503 -205 505 -200
rect 510 -205 512 -200
rect 517 -205 519 -200
rect 621 -197 623 -192
rect 557 -205 559 -200
rect 564 -205 566 -200
rect 571 -205 573 -200
rect 578 -205 580 -200
rect 588 -205 590 -200
rect 595 -205 597 -200
rect 602 -205 604 -200
rect 609 -205 611 -200
rect -679 -224 -677 -219
rect -653 -224 -651 -219
rect -631 -223 -629 -218
rect -521 -214 -519 -210
rect -514 -214 -512 -210
rect -486 -214 -484 -210
rect -479 -214 -477 -210
rect -619 -222 -617 -217
rect -609 -222 -607 -217
rect -599 -222 -597 -217
rect -679 -245 -677 -242
rect -653 -245 -651 -242
rect -631 -245 -629 -236
rect -619 -238 -617 -235
rect -623 -240 -617 -238
rect -623 -242 -621 -240
rect -619 -242 -617 -240
rect -623 -244 -617 -242
rect -683 -247 -677 -245
rect -683 -249 -681 -247
rect -679 -249 -677 -247
rect -683 -251 -677 -249
rect -657 -247 -651 -245
rect -657 -249 -655 -247
rect -653 -249 -651 -247
rect -657 -251 -651 -249
rect -635 -247 -629 -245
rect -635 -249 -633 -247
rect -631 -249 -629 -247
rect -635 -251 -624 -249
rect -679 -254 -677 -251
rect -653 -254 -651 -251
rect -626 -255 -624 -251
rect -619 -255 -617 -244
rect -609 -245 -607 -235
rect -577 -223 -575 -218
rect -565 -222 -563 -217
rect -555 -222 -553 -217
rect -545 -222 -543 -217
rect -599 -245 -597 -240
rect -577 -245 -575 -236
rect -565 -238 -563 -235
rect -569 -240 -563 -238
rect -569 -242 -567 -240
rect -565 -242 -563 -240
rect -569 -244 -563 -242
rect -613 -247 -607 -245
rect -613 -249 -611 -247
rect -609 -249 -607 -247
rect -613 -251 -607 -249
rect -603 -247 -597 -245
rect -603 -249 -601 -247
rect -599 -249 -597 -247
rect -603 -251 -597 -249
rect -581 -247 -575 -245
rect -581 -249 -579 -247
rect -577 -249 -575 -247
rect -581 -251 -570 -249
rect -612 -255 -610 -251
rect -599 -255 -597 -251
rect -572 -255 -570 -251
rect -565 -255 -563 -244
rect -555 -245 -553 -235
rect -545 -245 -543 -240
rect -451 -223 -449 -218
rect -439 -222 -437 -217
rect -429 -222 -427 -217
rect -419 -222 -417 -217
rect -559 -247 -553 -245
rect -559 -249 -557 -247
rect -555 -249 -553 -247
rect -559 -251 -553 -249
rect -549 -247 -543 -245
rect -549 -249 -547 -247
rect -545 -249 -543 -247
rect -521 -248 -519 -242
rect -514 -245 -512 -242
rect -549 -251 -543 -249
rect -558 -255 -556 -251
rect -545 -255 -543 -251
rect -525 -250 -519 -248
rect -525 -252 -523 -250
rect -521 -252 -519 -250
rect -515 -247 -509 -245
rect -515 -249 -513 -247
rect -511 -249 -509 -247
rect -486 -248 -484 -242
rect -479 -245 -477 -242
rect -451 -245 -449 -236
rect -439 -238 -437 -235
rect -443 -240 -437 -238
rect -443 -242 -441 -240
rect -439 -242 -437 -240
rect -443 -244 -437 -242
rect -515 -251 -509 -249
rect -490 -250 -484 -248
rect -525 -254 -519 -252
rect -679 -268 -677 -263
rect -653 -268 -651 -263
rect -626 -273 -624 -268
rect -619 -273 -617 -268
rect -612 -273 -610 -268
rect -599 -269 -597 -264
rect -523 -257 -521 -254
rect -572 -273 -570 -268
rect -565 -273 -563 -268
rect -558 -273 -556 -268
rect -545 -269 -543 -264
rect -512 -260 -510 -251
rect -490 -252 -488 -250
rect -486 -252 -484 -250
rect -480 -247 -474 -245
rect -480 -249 -478 -247
rect -476 -249 -474 -247
rect -480 -251 -474 -249
rect -455 -247 -449 -245
rect -455 -249 -453 -247
rect -451 -249 -449 -247
rect -455 -251 -444 -249
rect -490 -254 -484 -252
rect -488 -257 -486 -254
rect -523 -269 -521 -265
rect -477 -260 -475 -251
rect -446 -255 -444 -251
rect -439 -255 -437 -244
rect -429 -245 -427 -235
rect -394 -224 -392 -219
rect -419 -245 -417 -240
rect -368 -224 -366 -219
rect -346 -223 -344 -218
rect -236 -214 -234 -210
rect -229 -214 -227 -210
rect -201 -214 -199 -210
rect -194 -214 -192 -210
rect -334 -222 -332 -217
rect -324 -222 -322 -217
rect -314 -222 -312 -217
rect -394 -245 -392 -242
rect -368 -245 -366 -242
rect -346 -245 -344 -236
rect -334 -238 -332 -235
rect -338 -240 -332 -238
rect -338 -242 -336 -240
rect -334 -242 -332 -240
rect -338 -244 -332 -242
rect -433 -247 -427 -245
rect -433 -249 -431 -247
rect -429 -249 -427 -247
rect -433 -251 -427 -249
rect -423 -247 -417 -245
rect -423 -249 -421 -247
rect -419 -249 -417 -247
rect -423 -251 -417 -249
rect -398 -247 -392 -245
rect -398 -249 -396 -247
rect -394 -249 -392 -247
rect -398 -251 -392 -249
rect -372 -247 -366 -245
rect -372 -249 -370 -247
rect -368 -249 -366 -247
rect -372 -251 -366 -249
rect -350 -247 -344 -245
rect -350 -249 -348 -247
rect -346 -249 -344 -247
rect -350 -251 -339 -249
rect -432 -255 -430 -251
rect -419 -255 -417 -251
rect -394 -254 -392 -251
rect -368 -254 -366 -251
rect -512 -273 -510 -268
rect -488 -269 -486 -265
rect -341 -255 -339 -251
rect -334 -255 -332 -244
rect -324 -245 -322 -235
rect -292 -223 -290 -218
rect -280 -222 -278 -217
rect -270 -222 -268 -217
rect -260 -222 -258 -217
rect -314 -245 -312 -240
rect -292 -245 -290 -236
rect -280 -238 -278 -235
rect -284 -240 -278 -238
rect -284 -242 -282 -240
rect -280 -242 -278 -240
rect -284 -244 -278 -242
rect -328 -247 -322 -245
rect -328 -249 -326 -247
rect -324 -249 -322 -247
rect -328 -251 -322 -249
rect -318 -247 -312 -245
rect -318 -249 -316 -247
rect -314 -249 -312 -247
rect -318 -251 -312 -249
rect -296 -247 -290 -245
rect -296 -249 -294 -247
rect -292 -249 -290 -247
rect -296 -251 -285 -249
rect -327 -255 -325 -251
rect -314 -255 -312 -251
rect -287 -255 -285 -251
rect -280 -255 -278 -244
rect -270 -245 -268 -235
rect -260 -245 -258 -240
rect -166 -223 -164 -218
rect -154 -222 -152 -217
rect -144 -222 -142 -217
rect -134 -222 -132 -217
rect -274 -247 -268 -245
rect -274 -249 -272 -247
rect -270 -249 -268 -247
rect -274 -251 -268 -249
rect -264 -247 -258 -245
rect -264 -249 -262 -247
rect -260 -249 -258 -247
rect -236 -248 -234 -242
rect -229 -245 -227 -242
rect -264 -251 -258 -249
rect -273 -255 -271 -251
rect -260 -255 -258 -251
rect -240 -250 -234 -248
rect -240 -252 -238 -250
rect -236 -252 -234 -250
rect -230 -247 -224 -245
rect -230 -249 -228 -247
rect -226 -249 -224 -247
rect -201 -248 -199 -242
rect -194 -245 -192 -242
rect -166 -245 -164 -236
rect -154 -238 -152 -235
rect -158 -240 -152 -238
rect -158 -242 -156 -240
rect -154 -242 -152 -240
rect -158 -244 -152 -242
rect -230 -251 -224 -249
rect -205 -250 -199 -248
rect -240 -254 -234 -252
rect -477 -273 -475 -268
rect -446 -273 -444 -268
rect -439 -273 -437 -268
rect -432 -273 -430 -268
rect -419 -269 -417 -264
rect -394 -268 -392 -263
rect -368 -268 -366 -263
rect -341 -273 -339 -268
rect -334 -273 -332 -268
rect -327 -273 -325 -268
rect -314 -269 -312 -264
rect -238 -257 -236 -254
rect -287 -273 -285 -268
rect -280 -273 -278 -268
rect -273 -273 -271 -268
rect -260 -269 -258 -264
rect -227 -260 -225 -251
rect -205 -252 -203 -250
rect -201 -252 -199 -250
rect -195 -247 -189 -245
rect -195 -249 -193 -247
rect -191 -249 -189 -247
rect -195 -251 -189 -249
rect -170 -247 -164 -245
rect -170 -249 -168 -247
rect -166 -249 -164 -247
rect -170 -251 -159 -249
rect -205 -254 -199 -252
rect -203 -257 -201 -254
rect -238 -269 -236 -265
rect -192 -260 -190 -251
rect -161 -255 -159 -251
rect -154 -255 -152 -244
rect -144 -245 -142 -235
rect -109 -224 -107 -219
rect -134 -245 -132 -240
rect -83 -224 -81 -219
rect -61 -223 -59 -218
rect 49 -214 51 -210
rect 56 -214 58 -210
rect 84 -214 86 -210
rect 91 -214 93 -210
rect -49 -222 -47 -217
rect -39 -222 -37 -217
rect -29 -222 -27 -217
rect -109 -245 -107 -242
rect -83 -245 -81 -242
rect -61 -245 -59 -236
rect -49 -238 -47 -235
rect -53 -240 -47 -238
rect -53 -242 -51 -240
rect -49 -242 -47 -240
rect -53 -244 -47 -242
rect -148 -247 -142 -245
rect -148 -249 -146 -247
rect -144 -249 -142 -247
rect -148 -251 -142 -249
rect -138 -247 -132 -245
rect -138 -249 -136 -247
rect -134 -249 -132 -247
rect -138 -251 -132 -249
rect -113 -247 -107 -245
rect -113 -249 -111 -247
rect -109 -249 -107 -247
rect -113 -251 -107 -249
rect -87 -247 -81 -245
rect -87 -249 -85 -247
rect -83 -249 -81 -247
rect -87 -251 -81 -249
rect -65 -247 -59 -245
rect -65 -249 -63 -247
rect -61 -249 -59 -247
rect -65 -251 -54 -249
rect -147 -255 -145 -251
rect -134 -255 -132 -251
rect -109 -254 -107 -251
rect -83 -254 -81 -251
rect -227 -273 -225 -268
rect -203 -269 -201 -265
rect -56 -255 -54 -251
rect -49 -255 -47 -244
rect -39 -245 -37 -235
rect -7 -223 -5 -218
rect 5 -222 7 -217
rect 15 -222 17 -217
rect 25 -222 27 -217
rect -29 -245 -27 -240
rect -7 -245 -5 -236
rect 5 -238 7 -235
rect 1 -240 7 -238
rect 1 -242 3 -240
rect 5 -242 7 -240
rect 1 -244 7 -242
rect -43 -247 -37 -245
rect -43 -249 -41 -247
rect -39 -249 -37 -247
rect -43 -251 -37 -249
rect -33 -247 -27 -245
rect -33 -249 -31 -247
rect -29 -249 -27 -247
rect -33 -251 -27 -249
rect -11 -247 -5 -245
rect -11 -249 -9 -247
rect -7 -249 -5 -247
rect -11 -251 0 -249
rect -42 -255 -40 -251
rect -29 -255 -27 -251
rect -2 -255 0 -251
rect 5 -255 7 -244
rect 15 -245 17 -235
rect 25 -245 27 -240
rect 119 -223 121 -218
rect 131 -222 133 -217
rect 141 -222 143 -217
rect 151 -222 153 -217
rect 11 -247 17 -245
rect 11 -249 13 -247
rect 15 -249 17 -247
rect 11 -251 17 -249
rect 21 -247 27 -245
rect 21 -249 23 -247
rect 25 -249 27 -247
rect 49 -248 51 -242
rect 56 -245 58 -242
rect 21 -251 27 -249
rect 12 -255 14 -251
rect 25 -255 27 -251
rect 45 -250 51 -248
rect 45 -252 47 -250
rect 49 -252 51 -250
rect 55 -247 61 -245
rect 55 -249 57 -247
rect 59 -249 61 -247
rect 84 -248 86 -242
rect 91 -245 93 -242
rect 119 -245 121 -236
rect 131 -238 133 -235
rect 127 -240 133 -238
rect 127 -242 129 -240
rect 131 -242 133 -240
rect 127 -244 133 -242
rect 55 -251 61 -249
rect 80 -250 86 -248
rect 45 -254 51 -252
rect -192 -273 -190 -268
rect -161 -273 -159 -268
rect -154 -273 -152 -268
rect -147 -273 -145 -268
rect -134 -269 -132 -264
rect -109 -268 -107 -263
rect -83 -268 -81 -263
rect -56 -273 -54 -268
rect -49 -273 -47 -268
rect -42 -273 -40 -268
rect -29 -269 -27 -264
rect 47 -257 49 -254
rect -2 -273 0 -268
rect 5 -273 7 -268
rect 12 -273 14 -268
rect 25 -269 27 -264
rect 58 -260 60 -251
rect 80 -252 82 -250
rect 84 -252 86 -250
rect 90 -247 96 -245
rect 90 -249 92 -247
rect 94 -249 96 -247
rect 90 -251 96 -249
rect 115 -247 121 -245
rect 115 -249 117 -247
rect 119 -249 121 -247
rect 115 -251 126 -249
rect 80 -254 86 -252
rect 82 -257 84 -254
rect 47 -269 49 -265
rect 93 -260 95 -251
rect 124 -255 126 -251
rect 131 -255 133 -244
rect 141 -245 143 -235
rect 176 -224 178 -219
rect 151 -245 153 -240
rect 202 -224 204 -219
rect 224 -223 226 -218
rect 334 -214 336 -210
rect 341 -214 343 -210
rect 369 -214 371 -210
rect 376 -214 378 -210
rect 236 -222 238 -217
rect 246 -222 248 -217
rect 256 -222 258 -217
rect 176 -245 178 -242
rect 202 -245 204 -242
rect 224 -245 226 -236
rect 236 -238 238 -235
rect 232 -240 238 -238
rect 232 -242 234 -240
rect 236 -242 238 -240
rect 232 -244 238 -242
rect 137 -247 143 -245
rect 137 -249 139 -247
rect 141 -249 143 -247
rect 137 -251 143 -249
rect 147 -247 153 -245
rect 147 -249 149 -247
rect 151 -249 153 -247
rect 147 -251 153 -249
rect 172 -247 178 -245
rect 172 -249 174 -247
rect 176 -249 178 -247
rect 172 -251 178 -249
rect 198 -247 204 -245
rect 198 -249 200 -247
rect 202 -249 204 -247
rect 198 -251 204 -249
rect 220 -247 226 -245
rect 220 -249 222 -247
rect 224 -249 226 -247
rect 220 -251 231 -249
rect 138 -255 140 -251
rect 151 -255 153 -251
rect 176 -254 178 -251
rect 202 -254 204 -251
rect 58 -273 60 -268
rect 82 -269 84 -265
rect 229 -255 231 -251
rect 236 -255 238 -244
rect 246 -245 248 -235
rect 278 -223 280 -218
rect 290 -222 292 -217
rect 300 -222 302 -217
rect 310 -222 312 -217
rect 256 -245 258 -240
rect 278 -245 280 -236
rect 290 -238 292 -235
rect 286 -240 292 -238
rect 286 -242 288 -240
rect 290 -242 292 -240
rect 286 -244 292 -242
rect 242 -247 248 -245
rect 242 -249 244 -247
rect 246 -249 248 -247
rect 242 -251 248 -249
rect 252 -247 258 -245
rect 252 -249 254 -247
rect 256 -249 258 -247
rect 252 -251 258 -249
rect 274 -247 280 -245
rect 274 -249 276 -247
rect 278 -249 280 -247
rect 274 -251 285 -249
rect 243 -255 245 -251
rect 256 -255 258 -251
rect 283 -255 285 -251
rect 290 -255 292 -244
rect 300 -245 302 -235
rect 310 -245 312 -240
rect 404 -223 406 -218
rect 465 -216 467 -211
rect 472 -216 474 -211
rect 479 -216 481 -211
rect 486 -216 488 -211
rect 496 -216 498 -211
rect 503 -216 505 -211
rect 510 -216 512 -211
rect 517 -216 519 -211
rect 416 -222 418 -217
rect 426 -222 428 -217
rect 436 -222 438 -217
rect 296 -247 302 -245
rect 296 -249 298 -247
rect 300 -249 302 -247
rect 296 -251 302 -249
rect 306 -247 312 -245
rect 306 -249 308 -247
rect 310 -249 312 -247
rect 334 -248 336 -242
rect 341 -245 343 -242
rect 306 -251 312 -249
rect 297 -255 299 -251
rect 310 -255 312 -251
rect 330 -250 336 -248
rect 330 -252 332 -250
rect 334 -252 336 -250
rect 340 -247 346 -245
rect 340 -249 342 -247
rect 344 -249 346 -247
rect 369 -248 371 -242
rect 376 -245 378 -242
rect 404 -245 406 -236
rect 416 -238 418 -235
rect 412 -240 418 -238
rect 412 -242 414 -240
rect 416 -242 418 -240
rect 412 -244 418 -242
rect 340 -251 346 -249
rect 365 -250 371 -248
rect 330 -254 336 -252
rect 93 -273 95 -268
rect 124 -273 126 -268
rect 131 -273 133 -268
rect 138 -273 140 -268
rect 151 -269 153 -264
rect 176 -268 178 -263
rect 202 -268 204 -263
rect 229 -273 231 -268
rect 236 -273 238 -268
rect 243 -273 245 -268
rect 256 -269 258 -264
rect 332 -257 334 -254
rect 283 -273 285 -268
rect 290 -273 292 -268
rect 297 -273 299 -268
rect 310 -269 312 -264
rect 343 -260 345 -251
rect 365 -252 367 -250
rect 369 -252 371 -250
rect 375 -247 381 -245
rect 375 -249 377 -247
rect 379 -249 381 -247
rect 375 -251 381 -249
rect 400 -247 406 -245
rect 400 -249 402 -247
rect 404 -249 406 -247
rect 400 -251 411 -249
rect 365 -254 371 -252
rect 367 -257 369 -254
rect 332 -269 334 -265
rect 378 -260 380 -251
rect 409 -255 411 -251
rect 416 -255 418 -244
rect 426 -245 428 -235
rect 557 -216 559 -211
rect 564 -216 566 -211
rect 571 -216 573 -211
rect 578 -216 580 -211
rect 588 -216 590 -211
rect 595 -216 597 -211
rect 602 -216 604 -211
rect 609 -216 611 -211
rect 529 -224 531 -219
rect 465 -237 467 -234
rect 459 -239 467 -237
rect 436 -245 438 -240
rect 459 -241 461 -239
rect 463 -241 465 -239
rect 459 -243 465 -241
rect 472 -243 474 -234
rect 422 -247 428 -245
rect 422 -249 424 -247
rect 426 -249 428 -247
rect 422 -251 428 -249
rect 432 -247 438 -245
rect 432 -249 434 -247
rect 436 -249 438 -247
rect 469 -245 475 -243
rect 469 -247 471 -245
rect 473 -247 475 -245
rect 469 -249 475 -247
rect 432 -251 438 -249
rect 423 -255 425 -251
rect 436 -255 438 -251
rect 479 -253 481 -234
rect 486 -237 488 -234
rect 496 -237 498 -234
rect 475 -255 481 -253
rect 343 -273 345 -268
rect 367 -269 369 -265
rect 378 -273 380 -268
rect 409 -273 411 -268
rect 416 -273 418 -268
rect 423 -273 425 -268
rect 436 -269 438 -264
rect 475 -257 477 -255
rect 479 -257 481 -255
rect 475 -259 481 -257
rect 485 -239 498 -237
rect 485 -241 487 -239
rect 489 -241 491 -239
rect 485 -243 491 -241
rect 503 -243 505 -234
rect 485 -262 487 -243
rect 495 -245 505 -243
rect 495 -253 497 -245
rect 510 -249 512 -234
rect 517 -239 519 -234
rect 516 -241 522 -239
rect 516 -243 518 -241
rect 520 -243 522 -241
rect 621 -224 623 -219
rect 557 -237 559 -234
rect 551 -239 559 -237
rect 551 -241 553 -239
rect 555 -241 557 -239
rect 516 -245 522 -243
rect 491 -255 497 -253
rect 501 -251 512 -249
rect 501 -253 503 -251
rect 505 -253 509 -251
rect 501 -255 509 -253
rect 491 -257 493 -255
rect 495 -257 497 -255
rect 491 -259 497 -257
rect 495 -262 497 -259
rect 507 -262 509 -255
rect 517 -262 519 -245
rect 529 -250 531 -242
rect 551 -243 557 -241
rect 564 -243 566 -234
rect 561 -245 567 -243
rect 561 -247 563 -245
rect 565 -247 567 -245
rect 561 -249 567 -247
rect 525 -252 531 -250
rect 525 -254 527 -252
rect 529 -254 531 -252
rect 571 -253 573 -234
rect 578 -237 580 -234
rect 588 -237 590 -234
rect 525 -256 531 -254
rect 567 -255 573 -253
rect 529 -259 531 -256
rect 485 -273 487 -268
rect 495 -273 497 -268
rect 507 -273 509 -268
rect 517 -273 519 -268
rect 529 -273 531 -268
rect 567 -257 569 -255
rect 571 -257 573 -255
rect 567 -259 573 -257
rect 577 -239 590 -237
rect 577 -241 579 -239
rect 581 -241 583 -239
rect 577 -243 583 -241
rect 595 -243 597 -234
rect 577 -262 579 -243
rect 587 -245 597 -243
rect 587 -253 589 -245
rect 602 -249 604 -234
rect 609 -239 611 -234
rect 608 -241 614 -239
rect 608 -243 610 -241
rect 612 -243 614 -241
rect 608 -245 614 -243
rect 583 -255 589 -253
rect 593 -251 604 -249
rect 593 -253 595 -251
rect 597 -253 601 -251
rect 593 -255 601 -253
rect 583 -257 585 -255
rect 587 -257 589 -255
rect 583 -259 589 -257
rect 587 -262 589 -259
rect 599 -262 601 -255
rect 609 -262 611 -245
rect 621 -250 623 -242
rect 617 -252 623 -250
rect 617 -254 619 -252
rect 621 -254 623 -252
rect 617 -256 623 -254
rect 621 -259 623 -256
rect 577 -273 579 -268
rect 587 -273 589 -268
rect 599 -273 601 -268
rect 609 -273 611 -268
rect 621 -273 623 -268
<< ndif >>
rect -608 209 -601 211
rect -608 207 -605 209
rect -603 207 -601 209
rect -608 202 -601 207
rect -554 209 -547 211
rect -554 207 -551 209
rect -549 207 -547 209
rect -633 200 -626 202
rect -633 198 -631 200
rect -629 198 -626 200
rect -690 195 -679 197
rect -690 193 -688 195
rect -686 193 -679 195
rect -690 188 -679 193
rect -677 194 -672 197
rect -664 195 -653 197
rect -677 192 -670 194
rect -677 190 -674 192
rect -672 190 -670 192
rect -677 188 -670 190
rect -664 193 -662 195
rect -660 193 -653 195
rect -664 188 -653 193
rect -651 194 -646 197
rect -633 196 -626 198
rect -651 192 -644 194
rect -651 190 -648 192
rect -646 190 -644 192
rect -651 188 -644 190
rect -631 189 -626 196
rect -624 189 -619 202
rect -617 189 -612 202
rect -610 198 -601 202
rect -554 202 -547 207
rect -508 209 -502 211
rect -508 207 -506 209
rect -504 207 -502 209
rect -579 200 -572 202
rect -579 198 -577 200
rect -575 198 -572 200
rect -610 189 -599 198
rect -597 195 -592 198
rect -579 196 -572 198
rect -597 193 -590 195
rect -597 191 -594 193
rect -592 191 -590 193
rect -597 189 -590 191
rect -577 189 -572 196
rect -570 189 -565 202
rect -563 189 -558 202
rect -556 198 -547 202
rect -508 202 -502 207
rect -473 209 -467 211
rect -473 207 -471 209
rect -469 207 -467 209
rect -428 209 -421 211
rect -428 207 -425 209
rect -423 207 -421 209
rect -519 200 -512 202
rect -519 199 -517 200
rect -556 189 -545 198
rect -543 195 -538 198
rect -530 197 -523 199
rect -530 195 -528 197
rect -526 195 -523 197
rect -543 193 -536 195
rect -543 191 -540 193
rect -538 191 -536 193
rect -530 191 -523 195
rect -521 198 -517 199
rect -515 198 -512 200
rect -521 194 -512 198
rect -510 194 -502 202
rect -473 202 -467 207
rect -428 202 -421 207
rect -323 209 -316 211
rect -323 207 -320 209
rect -318 207 -316 209
rect -484 200 -477 202
rect -484 199 -482 200
rect -495 197 -488 199
rect -495 195 -493 197
rect -491 195 -488 197
rect -521 191 -516 194
rect -543 189 -536 191
rect -495 191 -488 195
rect -486 198 -482 199
rect -480 198 -477 200
rect -486 194 -477 198
rect -475 194 -467 202
rect -453 200 -446 202
rect -453 198 -451 200
rect -449 198 -446 200
rect -453 196 -446 198
rect -486 191 -481 194
rect -451 189 -446 196
rect -444 189 -439 202
rect -437 189 -432 202
rect -430 198 -421 202
rect -323 202 -316 207
rect -269 209 -262 211
rect -269 207 -266 209
rect -264 207 -262 209
rect -430 189 -419 198
rect -417 195 -412 198
rect -348 200 -341 202
rect -348 198 -346 200
rect -344 198 -341 200
rect -405 195 -394 197
rect -417 193 -410 195
rect -417 191 -414 193
rect -412 191 -410 193
rect -417 189 -410 191
rect -405 193 -403 195
rect -401 193 -394 195
rect -405 188 -394 193
rect -392 194 -387 197
rect -379 195 -368 197
rect -392 192 -385 194
rect -392 190 -389 192
rect -387 190 -385 192
rect -392 188 -385 190
rect -379 193 -377 195
rect -375 193 -368 195
rect -379 188 -368 193
rect -366 194 -361 197
rect -348 196 -341 198
rect -366 192 -359 194
rect -366 190 -363 192
rect -361 190 -359 192
rect -366 188 -359 190
rect -346 189 -341 196
rect -339 189 -334 202
rect -332 189 -327 202
rect -325 198 -316 202
rect -269 202 -262 207
rect -223 209 -217 211
rect -223 207 -221 209
rect -219 207 -217 209
rect -294 200 -287 202
rect -294 198 -292 200
rect -290 198 -287 200
rect -325 189 -314 198
rect -312 195 -307 198
rect -294 196 -287 198
rect -312 193 -305 195
rect -312 191 -309 193
rect -307 191 -305 193
rect -312 189 -305 191
rect -292 189 -287 196
rect -285 189 -280 202
rect -278 189 -273 202
rect -271 198 -262 202
rect -223 202 -217 207
rect -188 209 -182 211
rect -188 207 -186 209
rect -184 207 -182 209
rect -143 209 -136 211
rect -143 207 -140 209
rect -138 207 -136 209
rect -234 200 -227 202
rect -234 199 -232 200
rect -271 189 -260 198
rect -258 195 -253 198
rect -245 197 -238 199
rect -245 195 -243 197
rect -241 195 -238 197
rect -258 193 -251 195
rect -258 191 -255 193
rect -253 191 -251 193
rect -245 191 -238 195
rect -236 198 -232 199
rect -230 198 -227 200
rect -236 194 -227 198
rect -225 194 -217 202
rect -188 202 -182 207
rect -143 202 -136 207
rect -38 209 -31 211
rect -38 207 -35 209
rect -33 207 -31 209
rect -199 200 -192 202
rect -199 199 -197 200
rect -210 197 -203 199
rect -210 195 -208 197
rect -206 195 -203 197
rect -236 191 -231 194
rect -258 189 -251 191
rect -210 191 -203 195
rect -201 198 -197 199
rect -195 198 -192 200
rect -201 194 -192 198
rect -190 194 -182 202
rect -168 200 -161 202
rect -168 198 -166 200
rect -164 198 -161 200
rect -168 196 -161 198
rect -201 191 -196 194
rect -166 189 -161 196
rect -159 189 -154 202
rect -152 189 -147 202
rect -145 198 -136 202
rect -38 202 -31 207
rect 16 209 23 211
rect 16 207 19 209
rect 21 207 23 209
rect -145 189 -134 198
rect -132 195 -127 198
rect -63 200 -56 202
rect -63 198 -61 200
rect -59 198 -56 200
rect -120 195 -109 197
rect -132 193 -125 195
rect -132 191 -129 193
rect -127 191 -125 193
rect -132 189 -125 191
rect -120 193 -118 195
rect -116 193 -109 195
rect -120 188 -109 193
rect -107 194 -102 197
rect -94 195 -83 197
rect -107 192 -100 194
rect -107 190 -104 192
rect -102 190 -100 192
rect -107 188 -100 190
rect -94 193 -92 195
rect -90 193 -83 195
rect -94 188 -83 193
rect -81 194 -76 197
rect -63 196 -56 198
rect -81 192 -74 194
rect -81 190 -78 192
rect -76 190 -74 192
rect -81 188 -74 190
rect -61 189 -56 196
rect -54 189 -49 202
rect -47 189 -42 202
rect -40 198 -31 202
rect 16 202 23 207
rect 62 209 68 211
rect 62 207 64 209
rect 66 207 68 209
rect -9 200 -2 202
rect -9 198 -7 200
rect -5 198 -2 200
rect -40 189 -29 198
rect -27 195 -22 198
rect -9 196 -2 198
rect -27 193 -20 195
rect -27 191 -24 193
rect -22 191 -20 193
rect -27 189 -20 191
rect -7 189 -2 196
rect 0 189 5 202
rect 7 189 12 202
rect 14 198 23 202
rect 62 202 68 207
rect 97 209 103 211
rect 97 207 99 209
rect 101 207 103 209
rect 142 209 149 211
rect 142 207 145 209
rect 147 207 149 209
rect 51 200 58 202
rect 51 199 53 200
rect 14 189 25 198
rect 27 195 32 198
rect 40 197 47 199
rect 40 195 42 197
rect 44 195 47 197
rect 27 193 34 195
rect 27 191 30 193
rect 32 191 34 193
rect 40 191 47 195
rect 49 198 53 199
rect 55 198 58 200
rect 49 194 58 198
rect 60 194 68 202
rect 97 202 103 207
rect 142 202 149 207
rect 247 209 254 211
rect 247 207 250 209
rect 252 207 254 209
rect 86 200 93 202
rect 86 199 88 200
rect 75 197 82 199
rect 75 195 77 197
rect 79 195 82 197
rect 49 191 54 194
rect 27 189 34 191
rect 75 191 82 195
rect 84 198 88 199
rect 90 198 93 200
rect 84 194 93 198
rect 95 194 103 202
rect 117 200 124 202
rect 117 198 119 200
rect 121 198 124 200
rect 117 196 124 198
rect 84 191 89 194
rect 119 189 124 196
rect 126 189 131 202
rect 133 189 138 202
rect 140 198 149 202
rect 247 202 254 207
rect 301 209 308 211
rect 301 207 304 209
rect 306 207 308 209
rect 140 189 151 198
rect 153 195 158 198
rect 222 200 229 202
rect 222 198 224 200
rect 226 198 229 200
rect 165 195 176 197
rect 153 193 160 195
rect 153 191 156 193
rect 158 191 160 193
rect 153 189 160 191
rect 165 193 167 195
rect 169 193 176 195
rect 165 188 176 193
rect 178 194 183 197
rect 191 195 202 197
rect 178 192 185 194
rect 178 190 181 192
rect 183 190 185 192
rect 178 188 185 190
rect 191 193 193 195
rect 195 193 202 195
rect 191 188 202 193
rect 204 194 209 197
rect 222 196 229 198
rect 204 192 211 194
rect 204 190 207 192
rect 209 190 211 192
rect 204 188 211 190
rect 224 189 229 196
rect 231 189 236 202
rect 238 189 243 202
rect 245 198 254 202
rect 301 202 308 207
rect 347 209 353 211
rect 347 207 349 209
rect 351 207 353 209
rect 276 200 283 202
rect 276 198 278 200
rect 280 198 283 200
rect 245 189 256 198
rect 258 195 263 198
rect 276 196 283 198
rect 258 193 265 195
rect 258 191 261 193
rect 263 191 265 193
rect 258 189 265 191
rect 278 189 283 196
rect 285 189 290 202
rect 292 189 297 202
rect 299 198 308 202
rect 347 202 353 207
rect 382 209 388 211
rect 382 207 384 209
rect 386 207 388 209
rect 427 209 434 211
rect 427 207 430 209
rect 432 207 434 209
rect 336 200 343 202
rect 336 199 338 200
rect 299 189 310 198
rect 312 195 317 198
rect 325 197 332 199
rect 325 195 327 197
rect 329 195 332 197
rect 312 193 319 195
rect 312 191 315 193
rect 317 191 319 193
rect 325 191 332 195
rect 334 198 338 199
rect 340 198 343 200
rect 334 194 343 198
rect 345 194 353 202
rect 382 202 388 207
rect 427 202 434 207
rect 465 209 472 211
rect 465 207 467 209
rect 469 207 472 209
rect 371 200 378 202
rect 371 199 373 200
rect 360 197 367 199
rect 360 195 362 197
rect 364 195 367 197
rect 334 191 339 194
rect 312 189 319 191
rect 360 191 367 195
rect 369 198 373 199
rect 375 198 378 200
rect 369 194 378 198
rect 380 194 388 202
rect 402 200 409 202
rect 402 198 404 200
rect 406 198 409 200
rect 402 196 409 198
rect 369 191 374 194
rect 404 189 409 196
rect 411 189 416 202
rect 418 189 423 202
rect 425 198 434 202
rect 465 202 472 207
rect 525 209 532 211
rect 525 207 527 209
rect 529 207 532 209
rect 465 198 474 202
rect 425 189 436 198
rect 438 195 443 198
rect 456 195 461 198
rect 438 193 445 195
rect 438 191 441 193
rect 443 191 445 193
rect 438 189 445 191
rect 454 193 461 195
rect 454 191 456 193
rect 458 191 461 193
rect 454 189 461 191
rect 463 189 474 198
rect 476 189 481 202
rect 483 189 488 202
rect 490 200 497 202
rect 490 198 493 200
rect 495 198 497 200
rect 525 202 532 207
rect 525 198 534 202
rect 490 196 497 198
rect 490 189 495 196
rect 516 195 521 198
rect 514 193 521 195
rect 514 191 516 193
rect 518 191 521 193
rect 514 189 521 191
rect 523 189 534 198
rect 536 189 541 202
rect 543 189 548 202
rect 550 200 557 202
rect 550 198 553 200
rect 555 198 557 200
rect 550 196 557 198
rect 550 189 555 196
rect 582 194 587 197
rect 580 192 587 194
rect 580 190 582 192
rect 584 190 587 192
rect 580 188 587 190
rect 589 195 600 197
rect 589 193 596 195
rect 598 193 600 195
rect 589 188 600 193
rect -690 91 -679 96
rect -690 89 -688 91
rect -686 89 -679 91
rect -690 87 -679 89
rect -677 94 -670 96
rect -677 92 -674 94
rect -672 92 -670 94
rect -677 90 -670 92
rect -664 91 -653 96
rect -677 87 -672 90
rect -664 89 -662 91
rect -660 89 -653 91
rect -664 87 -653 89
rect -651 94 -644 96
rect -651 92 -648 94
rect -646 92 -644 94
rect -651 90 -644 92
rect -651 87 -646 90
rect -631 88 -626 95
rect -633 86 -626 88
rect -633 84 -631 86
rect -629 84 -626 86
rect -633 82 -626 84
rect -624 82 -619 95
rect -617 82 -612 95
rect -610 86 -599 95
rect -597 93 -590 95
rect -597 91 -594 93
rect -592 91 -590 93
rect -597 89 -590 91
rect -597 86 -592 89
rect -577 88 -572 95
rect -579 86 -572 88
rect -610 82 -601 86
rect -608 77 -601 82
rect -579 84 -577 86
rect -575 84 -572 86
rect -579 82 -572 84
rect -570 82 -565 95
rect -563 82 -558 95
rect -556 86 -545 95
rect -543 93 -536 95
rect -543 91 -540 93
rect -538 91 -536 93
rect -543 89 -536 91
rect -530 89 -523 93
rect -543 86 -538 89
rect -530 87 -528 89
rect -526 87 -523 89
rect -556 82 -547 86
rect -608 75 -605 77
rect -603 75 -601 77
rect -608 73 -601 75
rect -554 77 -547 82
rect -530 85 -523 87
rect -521 90 -516 93
rect -521 86 -512 90
rect -521 85 -517 86
rect -519 84 -517 85
rect -515 84 -512 86
rect -519 82 -512 84
rect -510 82 -502 90
rect -495 89 -488 93
rect -495 87 -493 89
rect -491 87 -488 89
rect -495 85 -488 87
rect -486 90 -481 93
rect -486 86 -477 90
rect -486 85 -482 86
rect -554 75 -551 77
rect -549 75 -547 77
rect -554 73 -547 75
rect -508 77 -502 82
rect -484 84 -482 85
rect -480 84 -477 86
rect -484 82 -477 84
rect -475 82 -467 90
rect -451 88 -446 95
rect -453 86 -446 88
rect -453 84 -451 86
rect -449 84 -446 86
rect -453 82 -446 84
rect -444 82 -439 95
rect -437 82 -432 95
rect -430 86 -419 95
rect -417 93 -410 95
rect -417 91 -414 93
rect -412 91 -410 93
rect -417 89 -410 91
rect -405 91 -394 96
rect -405 89 -403 91
rect -401 89 -394 91
rect -417 86 -412 89
rect -405 87 -394 89
rect -392 94 -385 96
rect -392 92 -389 94
rect -387 92 -385 94
rect -392 90 -385 92
rect -379 91 -368 96
rect -392 87 -387 90
rect -379 89 -377 91
rect -375 89 -368 91
rect -379 87 -368 89
rect -366 94 -359 96
rect -366 92 -363 94
rect -361 92 -359 94
rect -366 90 -359 92
rect -366 87 -361 90
rect -346 88 -341 95
rect -430 82 -421 86
rect -508 75 -506 77
rect -504 75 -502 77
rect -508 73 -502 75
rect -473 77 -467 82
rect -428 77 -421 82
rect -348 86 -341 88
rect -348 84 -346 86
rect -344 84 -341 86
rect -348 82 -341 84
rect -339 82 -334 95
rect -332 82 -327 95
rect -325 86 -314 95
rect -312 93 -305 95
rect -312 91 -309 93
rect -307 91 -305 93
rect -312 89 -305 91
rect -312 86 -307 89
rect -292 88 -287 95
rect -294 86 -287 88
rect -325 82 -316 86
rect -473 75 -471 77
rect -469 75 -467 77
rect -473 73 -467 75
rect -428 75 -425 77
rect -423 75 -421 77
rect -428 73 -421 75
rect -323 77 -316 82
rect -294 84 -292 86
rect -290 84 -287 86
rect -294 82 -287 84
rect -285 82 -280 95
rect -278 82 -273 95
rect -271 86 -260 95
rect -258 93 -251 95
rect -258 91 -255 93
rect -253 91 -251 93
rect -258 89 -251 91
rect -245 89 -238 93
rect -258 86 -253 89
rect -245 87 -243 89
rect -241 87 -238 89
rect -271 82 -262 86
rect -323 75 -320 77
rect -318 75 -316 77
rect -323 73 -316 75
rect -269 77 -262 82
rect -245 85 -238 87
rect -236 90 -231 93
rect -236 86 -227 90
rect -236 85 -232 86
rect -234 84 -232 85
rect -230 84 -227 86
rect -234 82 -227 84
rect -225 82 -217 90
rect -210 89 -203 93
rect -210 87 -208 89
rect -206 87 -203 89
rect -210 85 -203 87
rect -201 90 -196 93
rect -201 86 -192 90
rect -201 85 -197 86
rect -269 75 -266 77
rect -264 75 -262 77
rect -269 73 -262 75
rect -223 77 -217 82
rect -199 84 -197 85
rect -195 84 -192 86
rect -199 82 -192 84
rect -190 82 -182 90
rect -166 88 -161 95
rect -168 86 -161 88
rect -168 84 -166 86
rect -164 84 -161 86
rect -168 82 -161 84
rect -159 82 -154 95
rect -152 82 -147 95
rect -145 86 -134 95
rect -132 93 -125 95
rect -132 91 -129 93
rect -127 91 -125 93
rect -132 89 -125 91
rect -120 91 -109 96
rect -120 89 -118 91
rect -116 89 -109 91
rect -132 86 -127 89
rect -120 87 -109 89
rect -107 94 -100 96
rect -107 92 -104 94
rect -102 92 -100 94
rect -107 90 -100 92
rect -94 91 -83 96
rect -107 87 -102 90
rect -94 89 -92 91
rect -90 89 -83 91
rect -94 87 -83 89
rect -81 94 -74 96
rect -81 92 -78 94
rect -76 92 -74 94
rect -81 90 -74 92
rect -81 87 -76 90
rect -61 88 -56 95
rect -145 82 -136 86
rect -223 75 -221 77
rect -219 75 -217 77
rect -223 73 -217 75
rect -188 77 -182 82
rect -143 77 -136 82
rect -63 86 -56 88
rect -63 84 -61 86
rect -59 84 -56 86
rect -63 82 -56 84
rect -54 82 -49 95
rect -47 82 -42 95
rect -40 86 -29 95
rect -27 93 -20 95
rect -27 91 -24 93
rect -22 91 -20 93
rect -27 89 -20 91
rect -27 86 -22 89
rect -7 88 -2 95
rect -9 86 -2 88
rect -40 82 -31 86
rect -188 75 -186 77
rect -184 75 -182 77
rect -188 73 -182 75
rect -143 75 -140 77
rect -138 75 -136 77
rect -143 73 -136 75
rect -38 77 -31 82
rect -9 84 -7 86
rect -5 84 -2 86
rect -9 82 -2 84
rect 0 82 5 95
rect 7 82 12 95
rect 14 86 25 95
rect 27 93 34 95
rect 27 91 30 93
rect 32 91 34 93
rect 27 89 34 91
rect 40 89 47 93
rect 27 86 32 89
rect 40 87 42 89
rect 44 87 47 89
rect 14 82 23 86
rect -38 75 -35 77
rect -33 75 -31 77
rect -38 73 -31 75
rect 16 77 23 82
rect 40 85 47 87
rect 49 90 54 93
rect 49 86 58 90
rect 49 85 53 86
rect 51 84 53 85
rect 55 84 58 86
rect 51 82 58 84
rect 60 82 68 90
rect 75 89 82 93
rect 75 87 77 89
rect 79 87 82 89
rect 75 85 82 87
rect 84 90 89 93
rect 84 86 93 90
rect 84 85 88 86
rect 16 75 19 77
rect 21 75 23 77
rect 16 73 23 75
rect 62 77 68 82
rect 86 84 88 85
rect 90 84 93 86
rect 86 82 93 84
rect 95 82 103 90
rect 119 88 124 95
rect 117 86 124 88
rect 117 84 119 86
rect 121 84 124 86
rect 117 82 124 84
rect 126 82 131 95
rect 133 82 138 95
rect 140 86 151 95
rect 153 93 160 95
rect 153 91 156 93
rect 158 91 160 93
rect 153 89 160 91
rect 165 91 176 96
rect 165 89 167 91
rect 169 89 176 91
rect 153 86 158 89
rect 165 87 176 89
rect 178 94 185 96
rect 178 92 181 94
rect 183 92 185 94
rect 178 90 185 92
rect 191 91 202 96
rect 178 87 183 90
rect 191 89 193 91
rect 195 89 202 91
rect 191 87 202 89
rect 204 94 211 96
rect 204 92 207 94
rect 209 92 211 94
rect 204 90 211 92
rect 204 87 209 90
rect 224 88 229 95
rect 140 82 149 86
rect 62 75 64 77
rect 66 75 68 77
rect 62 73 68 75
rect 97 77 103 82
rect 142 77 149 82
rect 222 86 229 88
rect 222 84 224 86
rect 226 84 229 86
rect 222 82 229 84
rect 231 82 236 95
rect 238 82 243 95
rect 245 86 256 95
rect 258 93 265 95
rect 258 91 261 93
rect 263 91 265 93
rect 258 89 265 91
rect 258 86 263 89
rect 278 88 283 95
rect 276 86 283 88
rect 245 82 254 86
rect 97 75 99 77
rect 101 75 103 77
rect 97 73 103 75
rect 142 75 145 77
rect 147 75 149 77
rect 142 73 149 75
rect 247 77 254 82
rect 276 84 278 86
rect 280 84 283 86
rect 276 82 283 84
rect 285 82 290 95
rect 292 82 297 95
rect 299 86 310 95
rect 312 93 319 95
rect 312 91 315 93
rect 317 91 319 93
rect 312 89 319 91
rect 325 89 332 93
rect 312 86 317 89
rect 325 87 327 89
rect 329 87 332 89
rect 299 82 308 86
rect 247 75 250 77
rect 252 75 254 77
rect 247 73 254 75
rect 301 77 308 82
rect 325 85 332 87
rect 334 90 339 93
rect 334 86 343 90
rect 334 85 338 86
rect 336 84 338 85
rect 340 84 343 86
rect 336 82 343 84
rect 345 82 353 90
rect 360 89 367 93
rect 360 87 362 89
rect 364 87 367 89
rect 360 85 367 87
rect 369 90 374 93
rect 369 86 378 90
rect 369 85 373 86
rect 301 75 304 77
rect 306 75 308 77
rect 301 73 308 75
rect 347 77 353 82
rect 371 84 373 85
rect 375 84 378 86
rect 371 82 378 84
rect 380 82 388 90
rect 404 88 409 95
rect 402 86 409 88
rect 402 84 404 86
rect 406 84 409 86
rect 402 82 409 84
rect 411 82 416 95
rect 418 82 423 95
rect 425 86 436 95
rect 438 93 445 95
rect 438 91 441 93
rect 443 91 445 93
rect 438 89 445 91
rect 454 93 461 95
rect 454 91 456 93
rect 458 91 461 93
rect 454 89 461 91
rect 438 86 443 89
rect 456 86 461 89
rect 463 86 474 95
rect 425 82 434 86
rect 347 75 349 77
rect 351 75 353 77
rect 347 73 353 75
rect 382 77 388 82
rect 427 77 434 82
rect 465 82 474 86
rect 476 82 481 95
rect 483 82 488 95
rect 490 88 495 95
rect 514 93 521 95
rect 514 91 516 93
rect 518 91 521 93
rect 514 89 521 91
rect 490 86 497 88
rect 516 86 521 89
rect 523 86 534 95
rect 490 84 493 86
rect 495 84 497 86
rect 490 82 497 84
rect 382 75 384 77
rect 386 75 388 77
rect 382 73 388 75
rect 427 75 430 77
rect 432 75 434 77
rect 427 73 434 75
rect 465 77 472 82
rect 525 82 534 86
rect 536 82 541 95
rect 543 82 548 95
rect 550 88 555 95
rect 580 94 587 96
rect 580 92 582 94
rect 584 92 587 94
rect 580 90 587 92
rect 550 86 557 88
rect 582 87 587 90
rect 589 91 600 96
rect 589 89 596 91
rect 598 89 600 91
rect 589 87 600 89
rect 550 84 553 86
rect 555 84 557 86
rect 550 82 557 84
rect 465 75 467 77
rect 469 75 472 77
rect 465 73 472 75
rect 525 77 532 82
rect 525 75 527 77
rect 529 75 532 77
rect 525 73 532 75
rect -608 -141 -601 -139
rect -608 -143 -605 -141
rect -603 -143 -601 -141
rect -608 -148 -601 -143
rect -554 -141 -547 -139
rect -554 -143 -551 -141
rect -549 -143 -547 -141
rect -633 -150 -626 -148
rect -633 -152 -631 -150
rect -629 -152 -626 -150
rect -690 -155 -679 -153
rect -690 -157 -688 -155
rect -686 -157 -679 -155
rect -690 -162 -679 -157
rect -677 -156 -672 -153
rect -664 -155 -653 -153
rect -677 -158 -670 -156
rect -677 -160 -674 -158
rect -672 -160 -670 -158
rect -677 -162 -670 -160
rect -664 -157 -662 -155
rect -660 -157 -653 -155
rect -664 -162 -653 -157
rect -651 -156 -646 -153
rect -633 -154 -626 -152
rect -651 -158 -644 -156
rect -651 -160 -648 -158
rect -646 -160 -644 -158
rect -651 -162 -644 -160
rect -631 -161 -626 -154
rect -624 -161 -619 -148
rect -617 -161 -612 -148
rect -610 -152 -601 -148
rect -554 -148 -547 -143
rect -508 -141 -502 -139
rect -508 -143 -506 -141
rect -504 -143 -502 -141
rect -579 -150 -572 -148
rect -579 -152 -577 -150
rect -575 -152 -572 -150
rect -610 -161 -599 -152
rect -597 -155 -592 -152
rect -579 -154 -572 -152
rect -597 -157 -590 -155
rect -597 -159 -594 -157
rect -592 -159 -590 -157
rect -597 -161 -590 -159
rect -577 -161 -572 -154
rect -570 -161 -565 -148
rect -563 -161 -558 -148
rect -556 -152 -547 -148
rect -508 -148 -502 -143
rect -473 -141 -467 -139
rect -473 -143 -471 -141
rect -469 -143 -467 -141
rect -428 -141 -421 -139
rect -428 -143 -425 -141
rect -423 -143 -421 -141
rect -519 -150 -512 -148
rect -519 -151 -517 -150
rect -556 -161 -545 -152
rect -543 -155 -538 -152
rect -530 -153 -523 -151
rect -530 -155 -528 -153
rect -526 -155 -523 -153
rect -543 -157 -536 -155
rect -543 -159 -540 -157
rect -538 -159 -536 -157
rect -530 -159 -523 -155
rect -521 -152 -517 -151
rect -515 -152 -512 -150
rect -521 -156 -512 -152
rect -510 -156 -502 -148
rect -473 -148 -467 -143
rect -428 -148 -421 -143
rect -323 -141 -316 -139
rect -323 -143 -320 -141
rect -318 -143 -316 -141
rect -484 -150 -477 -148
rect -484 -151 -482 -150
rect -495 -153 -488 -151
rect -495 -155 -493 -153
rect -491 -155 -488 -153
rect -521 -159 -516 -156
rect -543 -161 -536 -159
rect -495 -159 -488 -155
rect -486 -152 -482 -151
rect -480 -152 -477 -150
rect -486 -156 -477 -152
rect -475 -156 -467 -148
rect -453 -150 -446 -148
rect -453 -152 -451 -150
rect -449 -152 -446 -150
rect -453 -154 -446 -152
rect -486 -159 -481 -156
rect -451 -161 -446 -154
rect -444 -161 -439 -148
rect -437 -161 -432 -148
rect -430 -152 -421 -148
rect -323 -148 -316 -143
rect -269 -141 -262 -139
rect -269 -143 -266 -141
rect -264 -143 -262 -141
rect -430 -161 -419 -152
rect -417 -155 -412 -152
rect -348 -150 -341 -148
rect -348 -152 -346 -150
rect -344 -152 -341 -150
rect -405 -155 -394 -153
rect -417 -157 -410 -155
rect -417 -159 -414 -157
rect -412 -159 -410 -157
rect -417 -161 -410 -159
rect -405 -157 -403 -155
rect -401 -157 -394 -155
rect -405 -162 -394 -157
rect -392 -156 -387 -153
rect -379 -155 -368 -153
rect -392 -158 -385 -156
rect -392 -160 -389 -158
rect -387 -160 -385 -158
rect -392 -162 -385 -160
rect -379 -157 -377 -155
rect -375 -157 -368 -155
rect -379 -162 -368 -157
rect -366 -156 -361 -153
rect -348 -154 -341 -152
rect -366 -158 -359 -156
rect -366 -160 -363 -158
rect -361 -160 -359 -158
rect -366 -162 -359 -160
rect -346 -161 -341 -154
rect -339 -161 -334 -148
rect -332 -161 -327 -148
rect -325 -152 -316 -148
rect -269 -148 -262 -143
rect -223 -141 -217 -139
rect -223 -143 -221 -141
rect -219 -143 -217 -141
rect -294 -150 -287 -148
rect -294 -152 -292 -150
rect -290 -152 -287 -150
rect -325 -161 -314 -152
rect -312 -155 -307 -152
rect -294 -154 -287 -152
rect -312 -157 -305 -155
rect -312 -159 -309 -157
rect -307 -159 -305 -157
rect -312 -161 -305 -159
rect -292 -161 -287 -154
rect -285 -161 -280 -148
rect -278 -161 -273 -148
rect -271 -152 -262 -148
rect -223 -148 -217 -143
rect -188 -141 -182 -139
rect -188 -143 -186 -141
rect -184 -143 -182 -141
rect -143 -141 -136 -139
rect -143 -143 -140 -141
rect -138 -143 -136 -141
rect -234 -150 -227 -148
rect -234 -151 -232 -150
rect -271 -161 -260 -152
rect -258 -155 -253 -152
rect -245 -153 -238 -151
rect -245 -155 -243 -153
rect -241 -155 -238 -153
rect -258 -157 -251 -155
rect -258 -159 -255 -157
rect -253 -159 -251 -157
rect -245 -159 -238 -155
rect -236 -152 -232 -151
rect -230 -152 -227 -150
rect -236 -156 -227 -152
rect -225 -156 -217 -148
rect -188 -148 -182 -143
rect -143 -148 -136 -143
rect -38 -141 -31 -139
rect -38 -143 -35 -141
rect -33 -143 -31 -141
rect -199 -150 -192 -148
rect -199 -151 -197 -150
rect -210 -153 -203 -151
rect -210 -155 -208 -153
rect -206 -155 -203 -153
rect -236 -159 -231 -156
rect -258 -161 -251 -159
rect -210 -159 -203 -155
rect -201 -152 -197 -151
rect -195 -152 -192 -150
rect -201 -156 -192 -152
rect -190 -156 -182 -148
rect -168 -150 -161 -148
rect -168 -152 -166 -150
rect -164 -152 -161 -150
rect -168 -154 -161 -152
rect -201 -159 -196 -156
rect -166 -161 -161 -154
rect -159 -161 -154 -148
rect -152 -161 -147 -148
rect -145 -152 -136 -148
rect -38 -148 -31 -143
rect 16 -141 23 -139
rect 16 -143 19 -141
rect 21 -143 23 -141
rect -145 -161 -134 -152
rect -132 -155 -127 -152
rect -63 -150 -56 -148
rect -63 -152 -61 -150
rect -59 -152 -56 -150
rect -120 -155 -109 -153
rect -132 -157 -125 -155
rect -132 -159 -129 -157
rect -127 -159 -125 -157
rect -132 -161 -125 -159
rect -120 -157 -118 -155
rect -116 -157 -109 -155
rect -120 -162 -109 -157
rect -107 -156 -102 -153
rect -94 -155 -83 -153
rect -107 -158 -100 -156
rect -107 -160 -104 -158
rect -102 -160 -100 -158
rect -107 -162 -100 -160
rect -94 -157 -92 -155
rect -90 -157 -83 -155
rect -94 -162 -83 -157
rect -81 -156 -76 -153
rect -63 -154 -56 -152
rect -81 -158 -74 -156
rect -81 -160 -78 -158
rect -76 -160 -74 -158
rect -81 -162 -74 -160
rect -61 -161 -56 -154
rect -54 -161 -49 -148
rect -47 -161 -42 -148
rect -40 -152 -31 -148
rect 16 -148 23 -143
rect 62 -141 68 -139
rect 62 -143 64 -141
rect 66 -143 68 -141
rect -9 -150 -2 -148
rect -9 -152 -7 -150
rect -5 -152 -2 -150
rect -40 -161 -29 -152
rect -27 -155 -22 -152
rect -9 -154 -2 -152
rect -27 -157 -20 -155
rect -27 -159 -24 -157
rect -22 -159 -20 -157
rect -27 -161 -20 -159
rect -7 -161 -2 -154
rect 0 -161 5 -148
rect 7 -161 12 -148
rect 14 -152 23 -148
rect 62 -148 68 -143
rect 97 -141 103 -139
rect 97 -143 99 -141
rect 101 -143 103 -141
rect 142 -141 149 -139
rect 142 -143 145 -141
rect 147 -143 149 -141
rect 51 -150 58 -148
rect 51 -151 53 -150
rect 14 -161 25 -152
rect 27 -155 32 -152
rect 40 -153 47 -151
rect 40 -155 42 -153
rect 44 -155 47 -153
rect 27 -157 34 -155
rect 27 -159 30 -157
rect 32 -159 34 -157
rect 40 -159 47 -155
rect 49 -152 53 -151
rect 55 -152 58 -150
rect 49 -156 58 -152
rect 60 -156 68 -148
rect 97 -148 103 -143
rect 142 -148 149 -143
rect 247 -141 254 -139
rect 247 -143 250 -141
rect 252 -143 254 -141
rect 86 -150 93 -148
rect 86 -151 88 -150
rect 75 -153 82 -151
rect 75 -155 77 -153
rect 79 -155 82 -153
rect 49 -159 54 -156
rect 27 -161 34 -159
rect 75 -159 82 -155
rect 84 -152 88 -151
rect 90 -152 93 -150
rect 84 -156 93 -152
rect 95 -156 103 -148
rect 117 -150 124 -148
rect 117 -152 119 -150
rect 121 -152 124 -150
rect 117 -154 124 -152
rect 84 -159 89 -156
rect 119 -161 124 -154
rect 126 -161 131 -148
rect 133 -161 138 -148
rect 140 -152 149 -148
rect 247 -148 254 -143
rect 301 -141 308 -139
rect 301 -143 304 -141
rect 306 -143 308 -141
rect 140 -161 151 -152
rect 153 -155 158 -152
rect 222 -150 229 -148
rect 222 -152 224 -150
rect 226 -152 229 -150
rect 165 -155 176 -153
rect 153 -157 160 -155
rect 153 -159 156 -157
rect 158 -159 160 -157
rect 153 -161 160 -159
rect 165 -157 167 -155
rect 169 -157 176 -155
rect 165 -162 176 -157
rect 178 -156 183 -153
rect 191 -155 202 -153
rect 178 -158 185 -156
rect 178 -160 181 -158
rect 183 -160 185 -158
rect 178 -162 185 -160
rect 191 -157 193 -155
rect 195 -157 202 -155
rect 191 -162 202 -157
rect 204 -156 209 -153
rect 222 -154 229 -152
rect 204 -158 211 -156
rect 204 -160 207 -158
rect 209 -160 211 -158
rect 204 -162 211 -160
rect 224 -161 229 -154
rect 231 -161 236 -148
rect 238 -161 243 -148
rect 245 -152 254 -148
rect 301 -148 308 -143
rect 347 -141 353 -139
rect 347 -143 349 -141
rect 351 -143 353 -141
rect 276 -150 283 -148
rect 276 -152 278 -150
rect 280 -152 283 -150
rect 245 -161 256 -152
rect 258 -155 263 -152
rect 276 -154 283 -152
rect 258 -157 265 -155
rect 258 -159 261 -157
rect 263 -159 265 -157
rect 258 -161 265 -159
rect 278 -161 283 -154
rect 285 -161 290 -148
rect 292 -161 297 -148
rect 299 -152 308 -148
rect 347 -148 353 -143
rect 382 -141 388 -139
rect 382 -143 384 -141
rect 386 -143 388 -141
rect 427 -141 434 -139
rect 427 -143 430 -141
rect 432 -143 434 -141
rect 336 -150 343 -148
rect 336 -151 338 -150
rect 299 -161 310 -152
rect 312 -155 317 -152
rect 325 -153 332 -151
rect 325 -155 327 -153
rect 329 -155 332 -153
rect 312 -157 319 -155
rect 312 -159 315 -157
rect 317 -159 319 -157
rect 325 -159 332 -155
rect 334 -152 338 -151
rect 340 -152 343 -150
rect 334 -156 343 -152
rect 345 -156 353 -148
rect 382 -148 388 -143
rect 427 -148 434 -143
rect 371 -150 378 -148
rect 371 -151 373 -150
rect 360 -153 367 -151
rect 360 -155 362 -153
rect 364 -155 367 -153
rect 334 -159 339 -156
rect 312 -161 319 -159
rect 360 -159 367 -155
rect 369 -152 373 -151
rect 375 -152 378 -150
rect 369 -156 378 -152
rect 380 -156 388 -148
rect 402 -150 409 -148
rect 402 -152 404 -150
rect 406 -152 409 -150
rect 402 -154 409 -152
rect 369 -159 374 -156
rect 404 -161 409 -154
rect 411 -161 416 -148
rect 418 -161 423 -148
rect 425 -152 434 -148
rect 425 -161 436 -152
rect 438 -155 443 -152
rect 438 -157 445 -155
rect 438 -159 441 -157
rect 443 -159 445 -157
rect 438 -161 445 -159
rect 477 -141 483 -139
rect 477 -143 479 -141
rect 481 -143 483 -141
rect 499 -141 505 -139
rect 499 -143 501 -141
rect 503 -143 505 -141
rect 521 -141 527 -139
rect 521 -143 523 -141
rect 525 -143 527 -141
rect 477 -148 483 -143
rect 499 -148 505 -143
rect 521 -148 527 -143
rect 477 -154 485 -148
rect 487 -150 495 -148
rect 487 -152 490 -150
rect 492 -152 495 -150
rect 487 -154 495 -152
rect 497 -154 507 -148
rect 509 -150 517 -148
rect 509 -152 512 -150
rect 514 -152 517 -150
rect 509 -154 517 -152
rect 519 -154 529 -148
rect 521 -157 529 -154
rect 531 -150 538 -148
rect 531 -152 534 -150
rect 536 -152 538 -150
rect 531 -154 538 -152
rect 531 -157 536 -154
rect 569 -141 575 -139
rect 569 -143 571 -141
rect 573 -143 575 -141
rect 591 -141 597 -139
rect 591 -143 593 -141
rect 595 -143 597 -141
rect 613 -141 619 -139
rect 613 -143 615 -141
rect 617 -143 619 -141
rect 569 -148 575 -143
rect 591 -148 597 -143
rect 613 -148 619 -143
rect 569 -154 577 -148
rect 579 -150 587 -148
rect 579 -152 582 -150
rect 584 -152 587 -150
rect 579 -154 587 -152
rect 589 -154 599 -148
rect 601 -150 609 -148
rect 601 -152 604 -150
rect 606 -152 609 -150
rect 601 -154 609 -152
rect 611 -154 621 -148
rect 613 -157 621 -154
rect 623 -150 630 -148
rect 623 -152 626 -150
rect 628 -152 630 -150
rect 623 -154 630 -152
rect 623 -157 628 -154
rect -690 -259 -679 -254
rect -690 -261 -688 -259
rect -686 -261 -679 -259
rect -690 -263 -679 -261
rect -677 -256 -670 -254
rect -677 -258 -674 -256
rect -672 -258 -670 -256
rect -677 -260 -670 -258
rect -664 -259 -653 -254
rect -677 -263 -672 -260
rect -664 -261 -662 -259
rect -660 -261 -653 -259
rect -664 -263 -653 -261
rect -651 -256 -644 -254
rect -651 -258 -648 -256
rect -646 -258 -644 -256
rect -651 -260 -644 -258
rect -651 -263 -646 -260
rect -631 -262 -626 -255
rect -633 -264 -626 -262
rect -633 -266 -631 -264
rect -629 -266 -626 -264
rect -633 -268 -626 -266
rect -624 -268 -619 -255
rect -617 -268 -612 -255
rect -610 -264 -599 -255
rect -597 -257 -590 -255
rect -597 -259 -594 -257
rect -592 -259 -590 -257
rect -597 -261 -590 -259
rect -597 -264 -592 -261
rect -577 -262 -572 -255
rect -579 -264 -572 -262
rect -610 -268 -601 -264
rect -608 -273 -601 -268
rect -579 -266 -577 -264
rect -575 -266 -572 -264
rect -579 -268 -572 -266
rect -570 -268 -565 -255
rect -563 -268 -558 -255
rect -556 -264 -545 -255
rect -543 -257 -536 -255
rect -543 -259 -540 -257
rect -538 -259 -536 -257
rect -543 -261 -536 -259
rect -530 -261 -523 -257
rect -543 -264 -538 -261
rect -530 -263 -528 -261
rect -526 -263 -523 -261
rect -556 -268 -547 -264
rect -608 -275 -605 -273
rect -603 -275 -601 -273
rect -608 -277 -601 -275
rect -554 -273 -547 -268
rect -530 -265 -523 -263
rect -521 -260 -516 -257
rect -521 -264 -512 -260
rect -521 -265 -517 -264
rect -519 -266 -517 -265
rect -515 -266 -512 -264
rect -519 -268 -512 -266
rect -510 -268 -502 -260
rect -495 -261 -488 -257
rect -495 -263 -493 -261
rect -491 -263 -488 -261
rect -495 -265 -488 -263
rect -486 -260 -481 -257
rect -486 -264 -477 -260
rect -486 -265 -482 -264
rect -554 -275 -551 -273
rect -549 -275 -547 -273
rect -554 -277 -547 -275
rect -508 -273 -502 -268
rect -484 -266 -482 -265
rect -480 -266 -477 -264
rect -484 -268 -477 -266
rect -475 -268 -467 -260
rect -451 -262 -446 -255
rect -453 -264 -446 -262
rect -453 -266 -451 -264
rect -449 -266 -446 -264
rect -453 -268 -446 -266
rect -444 -268 -439 -255
rect -437 -268 -432 -255
rect -430 -264 -419 -255
rect -417 -257 -410 -255
rect -417 -259 -414 -257
rect -412 -259 -410 -257
rect -417 -261 -410 -259
rect -405 -259 -394 -254
rect -405 -261 -403 -259
rect -401 -261 -394 -259
rect -417 -264 -412 -261
rect -405 -263 -394 -261
rect -392 -256 -385 -254
rect -392 -258 -389 -256
rect -387 -258 -385 -256
rect -392 -260 -385 -258
rect -379 -259 -368 -254
rect -392 -263 -387 -260
rect -379 -261 -377 -259
rect -375 -261 -368 -259
rect -379 -263 -368 -261
rect -366 -256 -359 -254
rect -366 -258 -363 -256
rect -361 -258 -359 -256
rect -366 -260 -359 -258
rect -366 -263 -361 -260
rect -346 -262 -341 -255
rect -430 -268 -421 -264
rect -508 -275 -506 -273
rect -504 -275 -502 -273
rect -508 -277 -502 -275
rect -473 -273 -467 -268
rect -428 -273 -421 -268
rect -348 -264 -341 -262
rect -348 -266 -346 -264
rect -344 -266 -341 -264
rect -348 -268 -341 -266
rect -339 -268 -334 -255
rect -332 -268 -327 -255
rect -325 -264 -314 -255
rect -312 -257 -305 -255
rect -312 -259 -309 -257
rect -307 -259 -305 -257
rect -312 -261 -305 -259
rect -312 -264 -307 -261
rect -292 -262 -287 -255
rect -294 -264 -287 -262
rect -325 -268 -316 -264
rect -473 -275 -471 -273
rect -469 -275 -467 -273
rect -473 -277 -467 -275
rect -428 -275 -425 -273
rect -423 -275 -421 -273
rect -428 -277 -421 -275
rect -323 -273 -316 -268
rect -294 -266 -292 -264
rect -290 -266 -287 -264
rect -294 -268 -287 -266
rect -285 -268 -280 -255
rect -278 -268 -273 -255
rect -271 -264 -260 -255
rect -258 -257 -251 -255
rect -258 -259 -255 -257
rect -253 -259 -251 -257
rect -258 -261 -251 -259
rect -245 -261 -238 -257
rect -258 -264 -253 -261
rect -245 -263 -243 -261
rect -241 -263 -238 -261
rect -271 -268 -262 -264
rect -323 -275 -320 -273
rect -318 -275 -316 -273
rect -323 -277 -316 -275
rect -269 -273 -262 -268
rect -245 -265 -238 -263
rect -236 -260 -231 -257
rect -236 -264 -227 -260
rect -236 -265 -232 -264
rect -234 -266 -232 -265
rect -230 -266 -227 -264
rect -234 -268 -227 -266
rect -225 -268 -217 -260
rect -210 -261 -203 -257
rect -210 -263 -208 -261
rect -206 -263 -203 -261
rect -210 -265 -203 -263
rect -201 -260 -196 -257
rect -201 -264 -192 -260
rect -201 -265 -197 -264
rect -269 -275 -266 -273
rect -264 -275 -262 -273
rect -269 -277 -262 -275
rect -223 -273 -217 -268
rect -199 -266 -197 -265
rect -195 -266 -192 -264
rect -199 -268 -192 -266
rect -190 -268 -182 -260
rect -166 -262 -161 -255
rect -168 -264 -161 -262
rect -168 -266 -166 -264
rect -164 -266 -161 -264
rect -168 -268 -161 -266
rect -159 -268 -154 -255
rect -152 -268 -147 -255
rect -145 -264 -134 -255
rect -132 -257 -125 -255
rect -132 -259 -129 -257
rect -127 -259 -125 -257
rect -132 -261 -125 -259
rect -120 -259 -109 -254
rect -120 -261 -118 -259
rect -116 -261 -109 -259
rect -132 -264 -127 -261
rect -120 -263 -109 -261
rect -107 -256 -100 -254
rect -107 -258 -104 -256
rect -102 -258 -100 -256
rect -107 -260 -100 -258
rect -94 -259 -83 -254
rect -107 -263 -102 -260
rect -94 -261 -92 -259
rect -90 -261 -83 -259
rect -94 -263 -83 -261
rect -81 -256 -74 -254
rect -81 -258 -78 -256
rect -76 -258 -74 -256
rect -81 -260 -74 -258
rect -81 -263 -76 -260
rect -61 -262 -56 -255
rect -145 -268 -136 -264
rect -223 -275 -221 -273
rect -219 -275 -217 -273
rect -223 -277 -217 -275
rect -188 -273 -182 -268
rect -143 -273 -136 -268
rect -63 -264 -56 -262
rect -63 -266 -61 -264
rect -59 -266 -56 -264
rect -63 -268 -56 -266
rect -54 -268 -49 -255
rect -47 -268 -42 -255
rect -40 -264 -29 -255
rect -27 -257 -20 -255
rect -27 -259 -24 -257
rect -22 -259 -20 -257
rect -27 -261 -20 -259
rect -27 -264 -22 -261
rect -7 -262 -2 -255
rect -9 -264 -2 -262
rect -40 -268 -31 -264
rect -188 -275 -186 -273
rect -184 -275 -182 -273
rect -188 -277 -182 -275
rect -143 -275 -140 -273
rect -138 -275 -136 -273
rect -143 -277 -136 -275
rect -38 -273 -31 -268
rect -9 -266 -7 -264
rect -5 -266 -2 -264
rect -9 -268 -2 -266
rect 0 -268 5 -255
rect 7 -268 12 -255
rect 14 -264 25 -255
rect 27 -257 34 -255
rect 27 -259 30 -257
rect 32 -259 34 -257
rect 27 -261 34 -259
rect 40 -261 47 -257
rect 27 -264 32 -261
rect 40 -263 42 -261
rect 44 -263 47 -261
rect 14 -268 23 -264
rect -38 -275 -35 -273
rect -33 -275 -31 -273
rect -38 -277 -31 -275
rect 16 -273 23 -268
rect 40 -265 47 -263
rect 49 -260 54 -257
rect 49 -264 58 -260
rect 49 -265 53 -264
rect 51 -266 53 -265
rect 55 -266 58 -264
rect 51 -268 58 -266
rect 60 -268 68 -260
rect 75 -261 82 -257
rect 75 -263 77 -261
rect 79 -263 82 -261
rect 75 -265 82 -263
rect 84 -260 89 -257
rect 84 -264 93 -260
rect 84 -265 88 -264
rect 16 -275 19 -273
rect 21 -275 23 -273
rect 16 -277 23 -275
rect 62 -273 68 -268
rect 86 -266 88 -265
rect 90 -266 93 -264
rect 86 -268 93 -266
rect 95 -268 103 -260
rect 119 -262 124 -255
rect 117 -264 124 -262
rect 117 -266 119 -264
rect 121 -266 124 -264
rect 117 -268 124 -266
rect 126 -268 131 -255
rect 133 -268 138 -255
rect 140 -264 151 -255
rect 153 -257 160 -255
rect 153 -259 156 -257
rect 158 -259 160 -257
rect 153 -261 160 -259
rect 165 -259 176 -254
rect 165 -261 167 -259
rect 169 -261 176 -259
rect 153 -264 158 -261
rect 165 -263 176 -261
rect 178 -256 185 -254
rect 178 -258 181 -256
rect 183 -258 185 -256
rect 178 -260 185 -258
rect 191 -259 202 -254
rect 178 -263 183 -260
rect 191 -261 193 -259
rect 195 -261 202 -259
rect 191 -263 202 -261
rect 204 -256 211 -254
rect 204 -258 207 -256
rect 209 -258 211 -256
rect 204 -260 211 -258
rect 204 -263 209 -260
rect 224 -262 229 -255
rect 140 -268 149 -264
rect 62 -275 64 -273
rect 66 -275 68 -273
rect 62 -277 68 -275
rect 97 -273 103 -268
rect 142 -273 149 -268
rect 222 -264 229 -262
rect 222 -266 224 -264
rect 226 -266 229 -264
rect 222 -268 229 -266
rect 231 -268 236 -255
rect 238 -268 243 -255
rect 245 -264 256 -255
rect 258 -257 265 -255
rect 258 -259 261 -257
rect 263 -259 265 -257
rect 258 -261 265 -259
rect 258 -264 263 -261
rect 278 -262 283 -255
rect 276 -264 283 -262
rect 245 -268 254 -264
rect 97 -275 99 -273
rect 101 -275 103 -273
rect 97 -277 103 -275
rect 142 -275 145 -273
rect 147 -275 149 -273
rect 142 -277 149 -275
rect 247 -273 254 -268
rect 276 -266 278 -264
rect 280 -266 283 -264
rect 276 -268 283 -266
rect 285 -268 290 -255
rect 292 -268 297 -255
rect 299 -264 310 -255
rect 312 -257 319 -255
rect 312 -259 315 -257
rect 317 -259 319 -257
rect 312 -261 319 -259
rect 325 -261 332 -257
rect 312 -264 317 -261
rect 325 -263 327 -261
rect 329 -263 332 -261
rect 299 -268 308 -264
rect 247 -275 250 -273
rect 252 -275 254 -273
rect 247 -277 254 -275
rect 301 -273 308 -268
rect 325 -265 332 -263
rect 334 -260 339 -257
rect 334 -264 343 -260
rect 334 -265 338 -264
rect 336 -266 338 -265
rect 340 -266 343 -264
rect 336 -268 343 -266
rect 345 -268 353 -260
rect 360 -261 367 -257
rect 360 -263 362 -261
rect 364 -263 367 -261
rect 360 -265 367 -263
rect 369 -260 374 -257
rect 369 -264 378 -260
rect 369 -265 373 -264
rect 301 -275 304 -273
rect 306 -275 308 -273
rect 301 -277 308 -275
rect 347 -273 353 -268
rect 371 -266 373 -265
rect 375 -266 378 -264
rect 371 -268 378 -266
rect 380 -268 388 -260
rect 404 -262 409 -255
rect 402 -264 409 -262
rect 402 -266 404 -264
rect 406 -266 409 -264
rect 402 -268 409 -266
rect 411 -268 416 -255
rect 418 -268 423 -255
rect 425 -264 436 -255
rect 438 -257 445 -255
rect 438 -259 441 -257
rect 443 -259 445 -257
rect 438 -261 445 -259
rect 438 -264 443 -261
rect 425 -268 434 -264
rect 347 -275 349 -273
rect 351 -275 353 -273
rect 347 -277 353 -275
rect 382 -273 388 -268
rect 427 -273 434 -268
rect 382 -275 384 -273
rect 386 -275 388 -273
rect 382 -277 388 -275
rect 427 -275 430 -273
rect 432 -275 434 -273
rect 427 -277 434 -275
rect 521 -262 529 -259
rect 477 -268 485 -262
rect 487 -264 495 -262
rect 487 -266 490 -264
rect 492 -266 495 -264
rect 487 -268 495 -266
rect 497 -268 507 -262
rect 509 -264 517 -262
rect 509 -266 512 -264
rect 514 -266 517 -264
rect 509 -268 517 -266
rect 519 -268 529 -262
rect 531 -262 536 -259
rect 531 -264 538 -262
rect 531 -266 534 -264
rect 536 -266 538 -264
rect 531 -268 538 -266
rect 477 -273 483 -268
rect 499 -273 505 -268
rect 521 -273 527 -268
rect 613 -262 621 -259
rect 477 -275 479 -273
rect 481 -275 483 -273
rect 477 -277 483 -275
rect 499 -275 501 -273
rect 503 -275 505 -273
rect 499 -277 505 -275
rect 521 -275 523 -273
rect 525 -275 527 -273
rect 521 -277 527 -275
rect 569 -268 577 -262
rect 579 -264 587 -262
rect 579 -266 582 -264
rect 584 -266 587 -264
rect 579 -268 587 -266
rect 589 -268 599 -262
rect 601 -264 609 -262
rect 601 -266 604 -264
rect 606 -266 609 -264
rect 601 -268 609 -266
rect 611 -268 621 -262
rect 623 -262 628 -259
rect 623 -264 630 -262
rect 623 -266 626 -264
rect 628 -266 630 -264
rect 623 -268 630 -266
rect 569 -273 575 -268
rect 591 -273 597 -268
rect 613 -273 619 -268
rect 569 -275 571 -273
rect 573 -275 575 -273
rect 569 -277 575 -275
rect 591 -275 593 -273
rect 595 -275 597 -273
rect 591 -277 597 -275
rect 613 -275 615 -273
rect 617 -275 619 -273
rect 613 -277 619 -275
<< pdif >>
rect -688 159 -679 176
rect -688 157 -685 159
rect -683 158 -679 159
rect -677 174 -670 176
rect -677 172 -674 174
rect -672 172 -670 174
rect -677 167 -670 172
rect -677 165 -674 167
rect -672 165 -670 167
rect -677 163 -670 165
rect -677 158 -672 163
rect -662 159 -653 176
rect -683 157 -681 158
rect -688 155 -681 157
rect -662 157 -659 159
rect -657 158 -653 159
rect -651 174 -644 176
rect -651 172 -648 174
rect -646 172 -644 174
rect -651 167 -644 172
rect -651 165 -648 167
rect -646 165 -644 167
rect -651 163 -644 165
rect -638 168 -631 170
rect -638 166 -636 168
rect -634 166 -631 168
rect -651 158 -646 163
rect -638 161 -631 166
rect -638 159 -636 161
rect -634 159 -631 161
rect -657 157 -655 158
rect -662 155 -655 157
rect -638 157 -631 159
rect -629 169 -624 170
rect -605 169 -599 174
rect -629 157 -619 169
rect -627 156 -619 157
rect -617 167 -609 169
rect -617 165 -614 167
rect -612 165 -609 167
rect -617 160 -609 165
rect -617 158 -614 160
rect -612 158 -609 160
rect -617 156 -609 158
rect -607 160 -599 169
rect -607 158 -604 160
rect -602 158 -599 160
rect -607 156 -599 158
rect -597 172 -590 174
rect -597 170 -594 172
rect -592 170 -590 172
rect -597 165 -590 170
rect -597 163 -594 165
rect -592 163 -590 165
rect -597 161 -590 163
rect -584 168 -577 170
rect -584 166 -582 168
rect -580 166 -577 168
rect -584 161 -577 166
rect -597 156 -592 161
rect -584 159 -582 161
rect -580 159 -577 161
rect -584 157 -577 159
rect -575 169 -570 170
rect -551 169 -545 174
rect -575 157 -565 169
rect -627 149 -621 156
rect -573 156 -565 157
rect -563 167 -555 169
rect -563 165 -560 167
rect -558 165 -555 167
rect -563 160 -555 165
rect -563 158 -560 160
rect -558 158 -555 160
rect -563 156 -555 158
rect -553 160 -545 169
rect -553 158 -550 160
rect -548 158 -545 160
rect -553 156 -545 158
rect -543 172 -536 174
rect -543 170 -540 172
rect -538 170 -536 172
rect -543 165 -536 170
rect -543 163 -540 165
rect -538 163 -536 165
rect -543 161 -536 163
rect -543 156 -538 161
rect -530 159 -521 176
rect -530 157 -528 159
rect -526 157 -521 159
rect -627 147 -625 149
rect -623 147 -621 149
rect -627 145 -621 147
rect -573 149 -567 156
rect -530 152 -521 157
rect -573 147 -571 149
rect -569 147 -567 149
rect -530 150 -528 152
rect -526 150 -521 152
rect -530 148 -521 150
rect -519 148 -514 176
rect -512 168 -507 176
rect -512 166 -505 168
rect -512 164 -509 166
rect -507 164 -505 166
rect -512 159 -505 164
rect -512 157 -509 159
rect -507 157 -505 159
rect -512 155 -505 157
rect -495 159 -486 176
rect -495 157 -493 159
rect -491 157 -486 159
rect -512 148 -507 155
rect -495 152 -486 157
rect -495 150 -493 152
rect -491 150 -486 152
rect -495 148 -486 150
rect -484 148 -479 176
rect -477 168 -472 176
rect -458 168 -451 170
rect -477 166 -470 168
rect -477 164 -474 166
rect -472 164 -470 166
rect -477 159 -470 164
rect -477 157 -474 159
rect -472 157 -470 159
rect -458 166 -456 168
rect -454 166 -451 168
rect -458 161 -451 166
rect -458 159 -456 161
rect -454 159 -451 161
rect -458 157 -451 159
rect -449 169 -444 170
rect -425 169 -419 174
rect -449 157 -439 169
rect -477 155 -470 157
rect -477 148 -472 155
rect -447 156 -439 157
rect -437 167 -429 169
rect -437 165 -434 167
rect -432 165 -429 167
rect -437 160 -429 165
rect -437 158 -434 160
rect -432 158 -429 160
rect -437 156 -429 158
rect -427 160 -419 169
rect -427 158 -424 160
rect -422 158 -419 160
rect -427 156 -419 158
rect -417 172 -410 174
rect -417 170 -414 172
rect -412 170 -410 172
rect -417 165 -410 170
rect -417 163 -414 165
rect -412 163 -410 165
rect -417 161 -410 163
rect -417 156 -412 161
rect -403 159 -394 176
rect -403 157 -400 159
rect -398 158 -394 159
rect -392 174 -385 176
rect -392 172 -389 174
rect -387 172 -385 174
rect -392 167 -385 172
rect -392 165 -389 167
rect -387 165 -385 167
rect -392 163 -385 165
rect -392 158 -387 163
rect -377 159 -368 176
rect -398 157 -396 158
rect -573 145 -567 147
rect -447 149 -441 156
rect -403 155 -396 157
rect -377 157 -374 159
rect -372 158 -368 159
rect -366 174 -359 176
rect -366 172 -363 174
rect -361 172 -359 174
rect -366 167 -359 172
rect -366 165 -363 167
rect -361 165 -359 167
rect -366 163 -359 165
rect -353 168 -346 170
rect -353 166 -351 168
rect -349 166 -346 168
rect -366 158 -361 163
rect -353 161 -346 166
rect -353 159 -351 161
rect -349 159 -346 161
rect -372 157 -370 158
rect -377 155 -370 157
rect -353 157 -346 159
rect -344 169 -339 170
rect -320 169 -314 174
rect -344 157 -334 169
rect -342 156 -334 157
rect -332 167 -324 169
rect -332 165 -329 167
rect -327 165 -324 167
rect -332 160 -324 165
rect -332 158 -329 160
rect -327 158 -324 160
rect -332 156 -324 158
rect -322 160 -314 169
rect -322 158 -319 160
rect -317 158 -314 160
rect -322 156 -314 158
rect -312 172 -305 174
rect -312 170 -309 172
rect -307 170 -305 172
rect -312 165 -305 170
rect -312 163 -309 165
rect -307 163 -305 165
rect -312 161 -305 163
rect -299 168 -292 170
rect -299 166 -297 168
rect -295 166 -292 168
rect -299 161 -292 166
rect -312 156 -307 161
rect -299 159 -297 161
rect -295 159 -292 161
rect -299 157 -292 159
rect -290 169 -285 170
rect -266 169 -260 174
rect -290 157 -280 169
rect -447 147 -445 149
rect -443 147 -441 149
rect -447 145 -441 147
rect -342 149 -336 156
rect -288 156 -280 157
rect -278 167 -270 169
rect -278 165 -275 167
rect -273 165 -270 167
rect -278 160 -270 165
rect -278 158 -275 160
rect -273 158 -270 160
rect -278 156 -270 158
rect -268 160 -260 169
rect -268 158 -265 160
rect -263 158 -260 160
rect -268 156 -260 158
rect -258 172 -251 174
rect -258 170 -255 172
rect -253 170 -251 172
rect -258 165 -251 170
rect -258 163 -255 165
rect -253 163 -251 165
rect -258 161 -251 163
rect -258 156 -253 161
rect -245 159 -236 176
rect -245 157 -243 159
rect -241 157 -236 159
rect -342 147 -340 149
rect -338 147 -336 149
rect -342 145 -336 147
rect -288 149 -282 156
rect -245 152 -236 157
rect -288 147 -286 149
rect -284 147 -282 149
rect -245 150 -243 152
rect -241 150 -236 152
rect -245 148 -236 150
rect -234 148 -229 176
rect -227 168 -222 176
rect -227 166 -220 168
rect -227 164 -224 166
rect -222 164 -220 166
rect -227 159 -220 164
rect -227 157 -224 159
rect -222 157 -220 159
rect -227 155 -220 157
rect -210 159 -201 176
rect -210 157 -208 159
rect -206 157 -201 159
rect -227 148 -222 155
rect -210 152 -201 157
rect -210 150 -208 152
rect -206 150 -201 152
rect -210 148 -201 150
rect -199 148 -194 176
rect -192 168 -187 176
rect -173 168 -166 170
rect -192 166 -185 168
rect -192 164 -189 166
rect -187 164 -185 166
rect -192 159 -185 164
rect -192 157 -189 159
rect -187 157 -185 159
rect -173 166 -171 168
rect -169 166 -166 168
rect -173 161 -166 166
rect -173 159 -171 161
rect -169 159 -166 161
rect -173 157 -166 159
rect -164 169 -159 170
rect -140 169 -134 174
rect -164 157 -154 169
rect -192 155 -185 157
rect -192 148 -187 155
rect -162 156 -154 157
rect -152 167 -144 169
rect -152 165 -149 167
rect -147 165 -144 167
rect -152 160 -144 165
rect -152 158 -149 160
rect -147 158 -144 160
rect -152 156 -144 158
rect -142 160 -134 169
rect -142 158 -139 160
rect -137 158 -134 160
rect -142 156 -134 158
rect -132 172 -125 174
rect -132 170 -129 172
rect -127 170 -125 172
rect -132 165 -125 170
rect -132 163 -129 165
rect -127 163 -125 165
rect -132 161 -125 163
rect -132 156 -127 161
rect -118 159 -109 176
rect -118 157 -115 159
rect -113 158 -109 159
rect -107 174 -100 176
rect -107 172 -104 174
rect -102 172 -100 174
rect -107 167 -100 172
rect -107 165 -104 167
rect -102 165 -100 167
rect -107 163 -100 165
rect -107 158 -102 163
rect -92 159 -83 176
rect -113 157 -111 158
rect -288 145 -282 147
rect -162 149 -156 156
rect -118 155 -111 157
rect -92 157 -89 159
rect -87 158 -83 159
rect -81 174 -74 176
rect -81 172 -78 174
rect -76 172 -74 174
rect -81 167 -74 172
rect -81 165 -78 167
rect -76 165 -74 167
rect -81 163 -74 165
rect -68 168 -61 170
rect -68 166 -66 168
rect -64 166 -61 168
rect -81 158 -76 163
rect -68 161 -61 166
rect -68 159 -66 161
rect -64 159 -61 161
rect -87 157 -85 158
rect -92 155 -85 157
rect -68 157 -61 159
rect -59 169 -54 170
rect -35 169 -29 174
rect -59 157 -49 169
rect -57 156 -49 157
rect -47 167 -39 169
rect -47 165 -44 167
rect -42 165 -39 167
rect -47 160 -39 165
rect -47 158 -44 160
rect -42 158 -39 160
rect -47 156 -39 158
rect -37 160 -29 169
rect -37 158 -34 160
rect -32 158 -29 160
rect -37 156 -29 158
rect -27 172 -20 174
rect -27 170 -24 172
rect -22 170 -20 172
rect -27 165 -20 170
rect -27 163 -24 165
rect -22 163 -20 165
rect -27 161 -20 163
rect -14 168 -7 170
rect -14 166 -12 168
rect -10 166 -7 168
rect -14 161 -7 166
rect -27 156 -22 161
rect -14 159 -12 161
rect -10 159 -7 161
rect -14 157 -7 159
rect -5 169 0 170
rect 19 169 25 174
rect -5 157 5 169
rect -162 147 -160 149
rect -158 147 -156 149
rect -162 145 -156 147
rect -57 149 -51 156
rect -3 156 5 157
rect 7 167 15 169
rect 7 165 10 167
rect 12 165 15 167
rect 7 160 15 165
rect 7 158 10 160
rect 12 158 15 160
rect 7 156 15 158
rect 17 160 25 169
rect 17 158 20 160
rect 22 158 25 160
rect 17 156 25 158
rect 27 172 34 174
rect 27 170 30 172
rect 32 170 34 172
rect 27 165 34 170
rect 27 163 30 165
rect 32 163 34 165
rect 27 161 34 163
rect 27 156 32 161
rect 40 159 49 176
rect 40 157 42 159
rect 44 157 49 159
rect -57 147 -55 149
rect -53 147 -51 149
rect -57 145 -51 147
rect -3 149 3 156
rect 40 152 49 157
rect -3 147 -1 149
rect 1 147 3 149
rect 40 150 42 152
rect 44 150 49 152
rect 40 148 49 150
rect 51 148 56 176
rect 58 168 63 176
rect 58 166 65 168
rect 58 164 61 166
rect 63 164 65 166
rect 58 159 65 164
rect 58 157 61 159
rect 63 157 65 159
rect 58 155 65 157
rect 75 159 84 176
rect 75 157 77 159
rect 79 157 84 159
rect 58 148 63 155
rect 75 152 84 157
rect 75 150 77 152
rect 79 150 84 152
rect 75 148 84 150
rect 86 148 91 176
rect 93 168 98 176
rect 112 168 119 170
rect 93 166 100 168
rect 93 164 96 166
rect 98 164 100 166
rect 93 159 100 164
rect 93 157 96 159
rect 98 157 100 159
rect 112 166 114 168
rect 116 166 119 168
rect 112 161 119 166
rect 112 159 114 161
rect 116 159 119 161
rect 112 157 119 159
rect 121 169 126 170
rect 145 169 151 174
rect 121 157 131 169
rect 93 155 100 157
rect 93 148 98 155
rect 123 156 131 157
rect 133 167 141 169
rect 133 165 136 167
rect 138 165 141 167
rect 133 160 141 165
rect 133 158 136 160
rect 138 158 141 160
rect 133 156 141 158
rect 143 160 151 169
rect 143 158 146 160
rect 148 158 151 160
rect 143 156 151 158
rect 153 172 160 174
rect 153 170 156 172
rect 158 170 160 172
rect 153 165 160 170
rect 153 163 156 165
rect 158 163 160 165
rect 153 161 160 163
rect 153 156 158 161
rect 167 159 176 176
rect 167 157 170 159
rect 172 158 176 159
rect 178 174 185 176
rect 178 172 181 174
rect 183 172 185 174
rect 178 167 185 172
rect 178 165 181 167
rect 183 165 185 167
rect 178 163 185 165
rect 178 158 183 163
rect 193 159 202 176
rect 172 157 174 158
rect -3 145 3 147
rect 123 149 129 156
rect 167 155 174 157
rect 193 157 196 159
rect 198 158 202 159
rect 204 174 211 176
rect 204 172 207 174
rect 209 172 211 174
rect 204 167 211 172
rect 204 165 207 167
rect 209 165 211 167
rect 204 163 211 165
rect 217 168 224 170
rect 217 166 219 168
rect 221 166 224 168
rect 204 158 209 163
rect 217 161 224 166
rect 217 159 219 161
rect 221 159 224 161
rect 198 157 200 158
rect 193 155 200 157
rect 217 157 224 159
rect 226 169 231 170
rect 250 169 256 174
rect 226 157 236 169
rect 228 156 236 157
rect 238 167 246 169
rect 238 165 241 167
rect 243 165 246 167
rect 238 160 246 165
rect 238 158 241 160
rect 243 158 246 160
rect 238 156 246 158
rect 248 160 256 169
rect 248 158 251 160
rect 253 158 256 160
rect 248 156 256 158
rect 258 172 265 174
rect 258 170 261 172
rect 263 170 265 172
rect 258 165 265 170
rect 258 163 261 165
rect 263 163 265 165
rect 258 161 265 163
rect 271 168 278 170
rect 271 166 273 168
rect 275 166 278 168
rect 271 161 278 166
rect 258 156 263 161
rect 271 159 273 161
rect 275 159 278 161
rect 271 157 278 159
rect 280 169 285 170
rect 304 169 310 174
rect 280 157 290 169
rect 123 147 125 149
rect 127 147 129 149
rect 123 145 129 147
rect 228 149 234 156
rect 282 156 290 157
rect 292 167 300 169
rect 292 165 295 167
rect 297 165 300 167
rect 292 160 300 165
rect 292 158 295 160
rect 297 158 300 160
rect 292 156 300 158
rect 302 160 310 169
rect 302 158 305 160
rect 307 158 310 160
rect 302 156 310 158
rect 312 172 319 174
rect 312 170 315 172
rect 317 170 319 172
rect 312 165 319 170
rect 312 163 315 165
rect 317 163 319 165
rect 312 161 319 163
rect 312 156 317 161
rect 325 159 334 176
rect 325 157 327 159
rect 329 157 334 159
rect 228 147 230 149
rect 232 147 234 149
rect 228 145 234 147
rect 282 149 288 156
rect 325 152 334 157
rect 282 147 284 149
rect 286 147 288 149
rect 325 150 327 152
rect 329 150 334 152
rect 325 148 334 150
rect 336 148 341 176
rect 343 168 348 176
rect 343 166 350 168
rect 343 164 346 166
rect 348 164 350 166
rect 343 159 350 164
rect 343 157 346 159
rect 348 157 350 159
rect 343 155 350 157
rect 360 159 369 176
rect 360 157 362 159
rect 364 157 369 159
rect 343 148 348 155
rect 360 152 369 157
rect 360 150 362 152
rect 364 150 369 152
rect 360 148 369 150
rect 371 148 376 176
rect 378 168 383 176
rect 397 168 404 170
rect 378 166 385 168
rect 378 164 381 166
rect 383 164 385 166
rect 378 159 385 164
rect 378 157 381 159
rect 383 157 385 159
rect 397 166 399 168
rect 401 166 404 168
rect 397 161 404 166
rect 397 159 399 161
rect 401 159 404 161
rect 397 157 404 159
rect 406 169 411 170
rect 430 169 436 174
rect 406 157 416 169
rect 378 155 385 157
rect 378 148 383 155
rect 408 156 416 157
rect 418 167 426 169
rect 418 165 421 167
rect 423 165 426 167
rect 418 160 426 165
rect 418 158 421 160
rect 423 158 426 160
rect 418 156 426 158
rect 428 160 436 169
rect 428 158 431 160
rect 433 158 436 160
rect 428 156 436 158
rect 438 172 445 174
rect 438 170 441 172
rect 443 170 445 172
rect 438 165 445 170
rect 438 163 441 165
rect 443 163 445 165
rect 438 161 445 163
rect 454 172 461 174
rect 454 170 456 172
rect 458 170 461 172
rect 454 165 461 170
rect 454 163 456 165
rect 458 163 461 165
rect 454 161 461 163
rect 438 156 443 161
rect 456 156 461 161
rect 463 169 469 174
rect 514 172 521 174
rect 514 170 516 172
rect 518 170 521 172
rect 488 169 493 170
rect 463 160 471 169
rect 463 158 466 160
rect 468 158 471 160
rect 463 156 471 158
rect 473 167 481 169
rect 473 165 476 167
rect 478 165 481 167
rect 473 160 481 165
rect 473 158 476 160
rect 478 158 481 160
rect 473 156 481 158
rect 483 157 493 169
rect 495 168 502 170
rect 495 166 498 168
rect 500 166 502 168
rect 495 161 502 166
rect 514 165 521 170
rect 514 163 516 165
rect 518 163 521 165
rect 514 161 521 163
rect 495 159 498 161
rect 500 159 502 161
rect 495 157 502 159
rect 483 156 491 157
rect 282 145 288 147
rect 408 149 414 156
rect 408 147 410 149
rect 412 147 414 149
rect 408 145 414 147
rect 485 149 491 156
rect 516 156 521 161
rect 523 169 529 174
rect 580 174 587 176
rect 580 172 582 174
rect 584 172 587 174
rect 548 169 553 170
rect 523 160 531 169
rect 523 158 526 160
rect 528 158 531 160
rect 523 156 531 158
rect 533 167 541 169
rect 533 165 536 167
rect 538 165 541 167
rect 533 160 541 165
rect 533 158 536 160
rect 538 158 541 160
rect 533 156 541 158
rect 543 157 553 169
rect 555 168 562 170
rect 555 166 558 168
rect 560 166 562 168
rect 555 161 562 166
rect 580 167 587 172
rect 580 165 582 167
rect 584 165 587 167
rect 580 163 587 165
rect 555 159 558 161
rect 560 159 562 161
rect 555 157 562 159
rect 582 158 587 163
rect 589 159 598 176
rect 589 158 593 159
rect 543 156 551 157
rect 485 147 487 149
rect 489 147 491 149
rect 485 145 491 147
rect 545 149 551 156
rect 591 157 593 158
rect 595 157 598 159
rect 591 155 598 157
rect 545 147 547 149
rect 549 147 551 149
rect 545 145 551 147
rect -627 137 -621 139
rect -627 135 -625 137
rect -623 135 -621 137
rect -688 127 -681 129
rect -688 125 -685 127
rect -683 126 -681 127
rect -662 127 -655 129
rect -683 125 -679 126
rect -688 108 -679 125
rect -677 121 -672 126
rect -662 125 -659 127
rect -657 126 -655 127
rect -627 128 -621 135
rect -573 137 -567 139
rect -573 135 -571 137
rect -569 135 -567 137
rect -627 127 -619 128
rect -657 125 -653 126
rect -677 119 -670 121
rect -677 117 -674 119
rect -672 117 -670 119
rect -677 112 -670 117
rect -677 110 -674 112
rect -672 110 -670 112
rect -677 108 -670 110
rect -662 108 -653 125
rect -651 121 -646 126
rect -638 125 -631 127
rect -638 123 -636 125
rect -634 123 -631 125
rect -651 119 -644 121
rect -651 117 -648 119
rect -646 117 -644 119
rect -651 112 -644 117
rect -638 118 -631 123
rect -638 116 -636 118
rect -634 116 -631 118
rect -638 114 -631 116
rect -629 115 -619 127
rect -617 126 -609 128
rect -617 124 -614 126
rect -612 124 -609 126
rect -617 119 -609 124
rect -617 117 -614 119
rect -612 117 -609 119
rect -617 115 -609 117
rect -607 126 -599 128
rect -607 124 -604 126
rect -602 124 -599 126
rect -607 115 -599 124
rect -629 114 -624 115
rect -651 110 -648 112
rect -646 110 -644 112
rect -651 108 -644 110
rect -605 110 -599 115
rect -597 123 -592 128
rect -573 128 -567 135
rect -530 134 -521 136
rect -530 132 -528 134
rect -526 132 -521 134
rect -573 127 -565 128
rect -584 125 -577 127
rect -584 123 -582 125
rect -580 123 -577 125
rect -597 121 -590 123
rect -597 119 -594 121
rect -592 119 -590 121
rect -597 114 -590 119
rect -584 118 -577 123
rect -584 116 -582 118
rect -580 116 -577 118
rect -584 114 -577 116
rect -575 115 -565 127
rect -563 126 -555 128
rect -563 124 -560 126
rect -558 124 -555 126
rect -563 119 -555 124
rect -563 117 -560 119
rect -558 117 -555 119
rect -563 115 -555 117
rect -553 126 -545 128
rect -553 124 -550 126
rect -548 124 -545 126
rect -553 115 -545 124
rect -575 114 -570 115
rect -597 112 -594 114
rect -592 112 -590 114
rect -597 110 -590 112
rect -551 110 -545 115
rect -543 123 -538 128
rect -530 127 -521 132
rect -530 125 -528 127
rect -526 125 -521 127
rect -543 121 -536 123
rect -543 119 -540 121
rect -538 119 -536 121
rect -543 114 -536 119
rect -543 112 -540 114
rect -538 112 -536 114
rect -543 110 -536 112
rect -530 108 -521 125
rect -519 108 -514 136
rect -512 129 -507 136
rect -495 134 -486 136
rect -495 132 -493 134
rect -491 132 -486 134
rect -512 127 -505 129
rect -512 125 -509 127
rect -507 125 -505 127
rect -512 120 -505 125
rect -512 118 -509 120
rect -507 118 -505 120
rect -512 116 -505 118
rect -495 127 -486 132
rect -495 125 -493 127
rect -491 125 -486 127
rect -512 108 -507 116
rect -495 108 -486 125
rect -484 108 -479 136
rect -477 129 -472 136
rect -447 137 -441 139
rect -447 135 -445 137
rect -443 135 -441 137
rect -477 127 -470 129
rect -447 128 -441 135
rect -342 137 -336 139
rect -342 135 -340 137
rect -338 135 -336 137
rect -447 127 -439 128
rect -477 125 -474 127
rect -472 125 -470 127
rect -477 120 -470 125
rect -477 118 -474 120
rect -472 118 -470 120
rect -477 116 -470 118
rect -458 125 -451 127
rect -458 123 -456 125
rect -454 123 -451 125
rect -458 118 -451 123
rect -458 116 -456 118
rect -454 116 -451 118
rect -477 108 -472 116
rect -458 114 -451 116
rect -449 115 -439 127
rect -437 126 -429 128
rect -437 124 -434 126
rect -432 124 -429 126
rect -437 119 -429 124
rect -437 117 -434 119
rect -432 117 -429 119
rect -437 115 -429 117
rect -427 126 -419 128
rect -427 124 -424 126
rect -422 124 -419 126
rect -427 115 -419 124
rect -449 114 -444 115
rect -425 110 -419 115
rect -417 123 -412 128
rect -403 127 -396 129
rect -403 125 -400 127
rect -398 126 -396 127
rect -377 127 -370 129
rect -398 125 -394 126
rect -417 121 -410 123
rect -417 119 -414 121
rect -412 119 -410 121
rect -417 114 -410 119
rect -417 112 -414 114
rect -412 112 -410 114
rect -417 110 -410 112
rect -403 108 -394 125
rect -392 121 -387 126
rect -377 125 -374 127
rect -372 126 -370 127
rect -342 128 -336 135
rect -288 137 -282 139
rect -288 135 -286 137
rect -284 135 -282 137
rect -342 127 -334 128
rect -372 125 -368 126
rect -392 119 -385 121
rect -392 117 -389 119
rect -387 117 -385 119
rect -392 112 -385 117
rect -392 110 -389 112
rect -387 110 -385 112
rect -392 108 -385 110
rect -377 108 -368 125
rect -366 121 -361 126
rect -353 125 -346 127
rect -353 123 -351 125
rect -349 123 -346 125
rect -366 119 -359 121
rect -366 117 -363 119
rect -361 117 -359 119
rect -366 112 -359 117
rect -353 118 -346 123
rect -353 116 -351 118
rect -349 116 -346 118
rect -353 114 -346 116
rect -344 115 -334 127
rect -332 126 -324 128
rect -332 124 -329 126
rect -327 124 -324 126
rect -332 119 -324 124
rect -332 117 -329 119
rect -327 117 -324 119
rect -332 115 -324 117
rect -322 126 -314 128
rect -322 124 -319 126
rect -317 124 -314 126
rect -322 115 -314 124
rect -344 114 -339 115
rect -366 110 -363 112
rect -361 110 -359 112
rect -366 108 -359 110
rect -320 110 -314 115
rect -312 123 -307 128
rect -288 128 -282 135
rect -245 134 -236 136
rect -245 132 -243 134
rect -241 132 -236 134
rect -288 127 -280 128
rect -299 125 -292 127
rect -299 123 -297 125
rect -295 123 -292 125
rect -312 121 -305 123
rect -312 119 -309 121
rect -307 119 -305 121
rect -312 114 -305 119
rect -299 118 -292 123
rect -299 116 -297 118
rect -295 116 -292 118
rect -299 114 -292 116
rect -290 115 -280 127
rect -278 126 -270 128
rect -278 124 -275 126
rect -273 124 -270 126
rect -278 119 -270 124
rect -278 117 -275 119
rect -273 117 -270 119
rect -278 115 -270 117
rect -268 126 -260 128
rect -268 124 -265 126
rect -263 124 -260 126
rect -268 115 -260 124
rect -290 114 -285 115
rect -312 112 -309 114
rect -307 112 -305 114
rect -312 110 -305 112
rect -266 110 -260 115
rect -258 123 -253 128
rect -245 127 -236 132
rect -245 125 -243 127
rect -241 125 -236 127
rect -258 121 -251 123
rect -258 119 -255 121
rect -253 119 -251 121
rect -258 114 -251 119
rect -258 112 -255 114
rect -253 112 -251 114
rect -258 110 -251 112
rect -245 108 -236 125
rect -234 108 -229 136
rect -227 129 -222 136
rect -210 134 -201 136
rect -210 132 -208 134
rect -206 132 -201 134
rect -227 127 -220 129
rect -227 125 -224 127
rect -222 125 -220 127
rect -227 120 -220 125
rect -227 118 -224 120
rect -222 118 -220 120
rect -227 116 -220 118
rect -210 127 -201 132
rect -210 125 -208 127
rect -206 125 -201 127
rect -227 108 -222 116
rect -210 108 -201 125
rect -199 108 -194 136
rect -192 129 -187 136
rect -162 137 -156 139
rect -162 135 -160 137
rect -158 135 -156 137
rect -192 127 -185 129
rect -162 128 -156 135
rect -57 137 -51 139
rect -57 135 -55 137
rect -53 135 -51 137
rect -162 127 -154 128
rect -192 125 -189 127
rect -187 125 -185 127
rect -192 120 -185 125
rect -192 118 -189 120
rect -187 118 -185 120
rect -192 116 -185 118
rect -173 125 -166 127
rect -173 123 -171 125
rect -169 123 -166 125
rect -173 118 -166 123
rect -173 116 -171 118
rect -169 116 -166 118
rect -192 108 -187 116
rect -173 114 -166 116
rect -164 115 -154 127
rect -152 126 -144 128
rect -152 124 -149 126
rect -147 124 -144 126
rect -152 119 -144 124
rect -152 117 -149 119
rect -147 117 -144 119
rect -152 115 -144 117
rect -142 126 -134 128
rect -142 124 -139 126
rect -137 124 -134 126
rect -142 115 -134 124
rect -164 114 -159 115
rect -140 110 -134 115
rect -132 123 -127 128
rect -118 127 -111 129
rect -118 125 -115 127
rect -113 126 -111 127
rect -92 127 -85 129
rect -113 125 -109 126
rect -132 121 -125 123
rect -132 119 -129 121
rect -127 119 -125 121
rect -132 114 -125 119
rect -132 112 -129 114
rect -127 112 -125 114
rect -132 110 -125 112
rect -118 108 -109 125
rect -107 121 -102 126
rect -92 125 -89 127
rect -87 126 -85 127
rect -57 128 -51 135
rect -3 137 3 139
rect -3 135 -1 137
rect 1 135 3 137
rect -57 127 -49 128
rect -87 125 -83 126
rect -107 119 -100 121
rect -107 117 -104 119
rect -102 117 -100 119
rect -107 112 -100 117
rect -107 110 -104 112
rect -102 110 -100 112
rect -107 108 -100 110
rect -92 108 -83 125
rect -81 121 -76 126
rect -68 125 -61 127
rect -68 123 -66 125
rect -64 123 -61 125
rect -81 119 -74 121
rect -81 117 -78 119
rect -76 117 -74 119
rect -81 112 -74 117
rect -68 118 -61 123
rect -68 116 -66 118
rect -64 116 -61 118
rect -68 114 -61 116
rect -59 115 -49 127
rect -47 126 -39 128
rect -47 124 -44 126
rect -42 124 -39 126
rect -47 119 -39 124
rect -47 117 -44 119
rect -42 117 -39 119
rect -47 115 -39 117
rect -37 126 -29 128
rect -37 124 -34 126
rect -32 124 -29 126
rect -37 115 -29 124
rect -59 114 -54 115
rect -81 110 -78 112
rect -76 110 -74 112
rect -81 108 -74 110
rect -35 110 -29 115
rect -27 123 -22 128
rect -3 128 3 135
rect 40 134 49 136
rect 40 132 42 134
rect 44 132 49 134
rect -3 127 5 128
rect -14 125 -7 127
rect -14 123 -12 125
rect -10 123 -7 125
rect -27 121 -20 123
rect -27 119 -24 121
rect -22 119 -20 121
rect -27 114 -20 119
rect -14 118 -7 123
rect -14 116 -12 118
rect -10 116 -7 118
rect -14 114 -7 116
rect -5 115 5 127
rect 7 126 15 128
rect 7 124 10 126
rect 12 124 15 126
rect 7 119 15 124
rect 7 117 10 119
rect 12 117 15 119
rect 7 115 15 117
rect 17 126 25 128
rect 17 124 20 126
rect 22 124 25 126
rect 17 115 25 124
rect -5 114 0 115
rect -27 112 -24 114
rect -22 112 -20 114
rect -27 110 -20 112
rect 19 110 25 115
rect 27 123 32 128
rect 40 127 49 132
rect 40 125 42 127
rect 44 125 49 127
rect 27 121 34 123
rect 27 119 30 121
rect 32 119 34 121
rect 27 114 34 119
rect 27 112 30 114
rect 32 112 34 114
rect 27 110 34 112
rect 40 108 49 125
rect 51 108 56 136
rect 58 129 63 136
rect 75 134 84 136
rect 75 132 77 134
rect 79 132 84 134
rect 58 127 65 129
rect 58 125 61 127
rect 63 125 65 127
rect 58 120 65 125
rect 58 118 61 120
rect 63 118 65 120
rect 58 116 65 118
rect 75 127 84 132
rect 75 125 77 127
rect 79 125 84 127
rect 58 108 63 116
rect 75 108 84 125
rect 86 108 91 136
rect 93 129 98 136
rect 123 137 129 139
rect 123 135 125 137
rect 127 135 129 137
rect 93 127 100 129
rect 123 128 129 135
rect 228 137 234 139
rect 228 135 230 137
rect 232 135 234 137
rect 123 127 131 128
rect 93 125 96 127
rect 98 125 100 127
rect 93 120 100 125
rect 93 118 96 120
rect 98 118 100 120
rect 93 116 100 118
rect 112 125 119 127
rect 112 123 114 125
rect 116 123 119 125
rect 112 118 119 123
rect 112 116 114 118
rect 116 116 119 118
rect 93 108 98 116
rect 112 114 119 116
rect 121 115 131 127
rect 133 126 141 128
rect 133 124 136 126
rect 138 124 141 126
rect 133 119 141 124
rect 133 117 136 119
rect 138 117 141 119
rect 133 115 141 117
rect 143 126 151 128
rect 143 124 146 126
rect 148 124 151 126
rect 143 115 151 124
rect 121 114 126 115
rect 145 110 151 115
rect 153 123 158 128
rect 167 127 174 129
rect 167 125 170 127
rect 172 126 174 127
rect 193 127 200 129
rect 172 125 176 126
rect 153 121 160 123
rect 153 119 156 121
rect 158 119 160 121
rect 153 114 160 119
rect 153 112 156 114
rect 158 112 160 114
rect 153 110 160 112
rect 167 108 176 125
rect 178 121 183 126
rect 193 125 196 127
rect 198 126 200 127
rect 228 128 234 135
rect 282 137 288 139
rect 282 135 284 137
rect 286 135 288 137
rect 228 127 236 128
rect 198 125 202 126
rect 178 119 185 121
rect 178 117 181 119
rect 183 117 185 119
rect 178 112 185 117
rect 178 110 181 112
rect 183 110 185 112
rect 178 108 185 110
rect 193 108 202 125
rect 204 121 209 126
rect 217 125 224 127
rect 217 123 219 125
rect 221 123 224 125
rect 204 119 211 121
rect 204 117 207 119
rect 209 117 211 119
rect 204 112 211 117
rect 217 118 224 123
rect 217 116 219 118
rect 221 116 224 118
rect 217 114 224 116
rect 226 115 236 127
rect 238 126 246 128
rect 238 124 241 126
rect 243 124 246 126
rect 238 119 246 124
rect 238 117 241 119
rect 243 117 246 119
rect 238 115 246 117
rect 248 126 256 128
rect 248 124 251 126
rect 253 124 256 126
rect 248 115 256 124
rect 226 114 231 115
rect 204 110 207 112
rect 209 110 211 112
rect 204 108 211 110
rect 250 110 256 115
rect 258 123 263 128
rect 282 128 288 135
rect 325 134 334 136
rect 325 132 327 134
rect 329 132 334 134
rect 282 127 290 128
rect 271 125 278 127
rect 271 123 273 125
rect 275 123 278 125
rect 258 121 265 123
rect 258 119 261 121
rect 263 119 265 121
rect 258 114 265 119
rect 271 118 278 123
rect 271 116 273 118
rect 275 116 278 118
rect 271 114 278 116
rect 280 115 290 127
rect 292 126 300 128
rect 292 124 295 126
rect 297 124 300 126
rect 292 119 300 124
rect 292 117 295 119
rect 297 117 300 119
rect 292 115 300 117
rect 302 126 310 128
rect 302 124 305 126
rect 307 124 310 126
rect 302 115 310 124
rect 280 114 285 115
rect 258 112 261 114
rect 263 112 265 114
rect 258 110 265 112
rect 304 110 310 115
rect 312 123 317 128
rect 325 127 334 132
rect 325 125 327 127
rect 329 125 334 127
rect 312 121 319 123
rect 312 119 315 121
rect 317 119 319 121
rect 312 114 319 119
rect 312 112 315 114
rect 317 112 319 114
rect 312 110 319 112
rect 325 108 334 125
rect 336 108 341 136
rect 343 129 348 136
rect 360 134 369 136
rect 360 132 362 134
rect 364 132 369 134
rect 343 127 350 129
rect 343 125 346 127
rect 348 125 350 127
rect 343 120 350 125
rect 343 118 346 120
rect 348 118 350 120
rect 343 116 350 118
rect 360 127 369 132
rect 360 125 362 127
rect 364 125 369 127
rect 343 108 348 116
rect 360 108 369 125
rect 371 108 376 136
rect 378 129 383 136
rect 408 137 414 139
rect 408 135 410 137
rect 412 135 414 137
rect 378 127 385 129
rect 408 128 414 135
rect 485 137 491 139
rect 485 135 487 137
rect 489 135 491 137
rect 485 128 491 135
rect 545 137 551 139
rect 545 135 547 137
rect 549 135 551 137
rect 408 127 416 128
rect 378 125 381 127
rect 383 125 385 127
rect 378 120 385 125
rect 378 118 381 120
rect 383 118 385 120
rect 378 116 385 118
rect 397 125 404 127
rect 397 123 399 125
rect 401 123 404 125
rect 397 118 404 123
rect 397 116 399 118
rect 401 116 404 118
rect 378 108 383 116
rect 397 114 404 116
rect 406 115 416 127
rect 418 126 426 128
rect 418 124 421 126
rect 423 124 426 126
rect 418 119 426 124
rect 418 117 421 119
rect 423 117 426 119
rect 418 115 426 117
rect 428 126 436 128
rect 428 124 431 126
rect 433 124 436 126
rect 428 115 436 124
rect 406 114 411 115
rect 430 110 436 115
rect 438 123 443 128
rect 456 123 461 128
rect 438 121 445 123
rect 438 119 441 121
rect 443 119 445 121
rect 438 114 445 119
rect 438 112 441 114
rect 443 112 445 114
rect 438 110 445 112
rect 454 121 461 123
rect 454 119 456 121
rect 458 119 461 121
rect 454 114 461 119
rect 454 112 456 114
rect 458 112 461 114
rect 454 110 461 112
rect 463 126 471 128
rect 463 124 466 126
rect 468 124 471 126
rect 463 115 471 124
rect 473 126 481 128
rect 473 124 476 126
rect 478 124 481 126
rect 473 119 481 124
rect 473 117 476 119
rect 478 117 481 119
rect 473 115 481 117
rect 483 127 491 128
rect 545 128 551 135
rect 483 115 493 127
rect 463 110 469 115
rect 488 114 493 115
rect 495 125 502 127
rect 495 123 498 125
rect 500 123 502 125
rect 516 123 521 128
rect 495 118 502 123
rect 495 116 498 118
rect 500 116 502 118
rect 495 114 502 116
rect 514 121 521 123
rect 514 119 516 121
rect 518 119 521 121
rect 514 114 521 119
rect 514 112 516 114
rect 518 112 521 114
rect 514 110 521 112
rect 523 126 531 128
rect 523 124 526 126
rect 528 124 531 126
rect 523 115 531 124
rect 533 126 541 128
rect 533 124 536 126
rect 538 124 541 126
rect 533 119 541 124
rect 533 117 536 119
rect 538 117 541 119
rect 533 115 541 117
rect 543 127 551 128
rect 543 115 553 127
rect 523 110 529 115
rect 548 114 553 115
rect 555 125 562 127
rect 591 127 598 129
rect 591 126 593 127
rect 555 123 558 125
rect 560 123 562 125
rect 555 118 562 123
rect 582 121 587 126
rect 555 116 558 118
rect 560 116 562 118
rect 555 114 562 116
rect 580 119 587 121
rect 580 117 582 119
rect 584 117 587 119
rect 580 112 587 117
rect 580 110 582 112
rect 584 110 587 112
rect 580 108 587 110
rect 589 125 593 126
rect 595 125 598 127
rect 589 108 598 125
rect -688 -191 -679 -174
rect -688 -193 -685 -191
rect -683 -192 -679 -191
rect -677 -176 -670 -174
rect -677 -178 -674 -176
rect -672 -178 -670 -176
rect -677 -183 -670 -178
rect -677 -185 -674 -183
rect -672 -185 -670 -183
rect -677 -187 -670 -185
rect -677 -192 -672 -187
rect -662 -191 -653 -174
rect -683 -193 -681 -192
rect -688 -195 -681 -193
rect -662 -193 -659 -191
rect -657 -192 -653 -191
rect -651 -176 -644 -174
rect -651 -178 -648 -176
rect -646 -178 -644 -176
rect -651 -183 -644 -178
rect -651 -185 -648 -183
rect -646 -185 -644 -183
rect -651 -187 -644 -185
rect -638 -182 -631 -180
rect -638 -184 -636 -182
rect -634 -184 -631 -182
rect -651 -192 -646 -187
rect -638 -189 -631 -184
rect -638 -191 -636 -189
rect -634 -191 -631 -189
rect -657 -193 -655 -192
rect -662 -195 -655 -193
rect -638 -193 -631 -191
rect -629 -181 -624 -180
rect -605 -181 -599 -176
rect -629 -193 -619 -181
rect -627 -194 -619 -193
rect -617 -183 -609 -181
rect -617 -185 -614 -183
rect -612 -185 -609 -183
rect -617 -190 -609 -185
rect -617 -192 -614 -190
rect -612 -192 -609 -190
rect -617 -194 -609 -192
rect -607 -190 -599 -181
rect -607 -192 -604 -190
rect -602 -192 -599 -190
rect -607 -194 -599 -192
rect -597 -178 -590 -176
rect -597 -180 -594 -178
rect -592 -180 -590 -178
rect -597 -185 -590 -180
rect -597 -187 -594 -185
rect -592 -187 -590 -185
rect -597 -189 -590 -187
rect -584 -182 -577 -180
rect -584 -184 -582 -182
rect -580 -184 -577 -182
rect -584 -189 -577 -184
rect -597 -194 -592 -189
rect -584 -191 -582 -189
rect -580 -191 -577 -189
rect -584 -193 -577 -191
rect -575 -181 -570 -180
rect -551 -181 -545 -176
rect -575 -193 -565 -181
rect -627 -201 -621 -194
rect -573 -194 -565 -193
rect -563 -183 -555 -181
rect -563 -185 -560 -183
rect -558 -185 -555 -183
rect -563 -190 -555 -185
rect -563 -192 -560 -190
rect -558 -192 -555 -190
rect -563 -194 -555 -192
rect -553 -190 -545 -181
rect -553 -192 -550 -190
rect -548 -192 -545 -190
rect -553 -194 -545 -192
rect -543 -178 -536 -176
rect -543 -180 -540 -178
rect -538 -180 -536 -178
rect -543 -185 -536 -180
rect -543 -187 -540 -185
rect -538 -187 -536 -185
rect -543 -189 -536 -187
rect -543 -194 -538 -189
rect -530 -191 -521 -174
rect -530 -193 -528 -191
rect -526 -193 -521 -191
rect -627 -203 -625 -201
rect -623 -203 -621 -201
rect -627 -205 -621 -203
rect -573 -201 -567 -194
rect -530 -198 -521 -193
rect -573 -203 -571 -201
rect -569 -203 -567 -201
rect -530 -200 -528 -198
rect -526 -200 -521 -198
rect -530 -202 -521 -200
rect -519 -202 -514 -174
rect -512 -182 -507 -174
rect -512 -184 -505 -182
rect -512 -186 -509 -184
rect -507 -186 -505 -184
rect -512 -191 -505 -186
rect -512 -193 -509 -191
rect -507 -193 -505 -191
rect -512 -195 -505 -193
rect -495 -191 -486 -174
rect -495 -193 -493 -191
rect -491 -193 -486 -191
rect -512 -202 -507 -195
rect -495 -198 -486 -193
rect -495 -200 -493 -198
rect -491 -200 -486 -198
rect -495 -202 -486 -200
rect -484 -202 -479 -174
rect -477 -182 -472 -174
rect -458 -182 -451 -180
rect -477 -184 -470 -182
rect -477 -186 -474 -184
rect -472 -186 -470 -184
rect -477 -191 -470 -186
rect -477 -193 -474 -191
rect -472 -193 -470 -191
rect -458 -184 -456 -182
rect -454 -184 -451 -182
rect -458 -189 -451 -184
rect -458 -191 -456 -189
rect -454 -191 -451 -189
rect -458 -193 -451 -191
rect -449 -181 -444 -180
rect -425 -181 -419 -176
rect -449 -193 -439 -181
rect -477 -195 -470 -193
rect -477 -202 -472 -195
rect -447 -194 -439 -193
rect -437 -183 -429 -181
rect -437 -185 -434 -183
rect -432 -185 -429 -183
rect -437 -190 -429 -185
rect -437 -192 -434 -190
rect -432 -192 -429 -190
rect -437 -194 -429 -192
rect -427 -190 -419 -181
rect -427 -192 -424 -190
rect -422 -192 -419 -190
rect -427 -194 -419 -192
rect -417 -178 -410 -176
rect -417 -180 -414 -178
rect -412 -180 -410 -178
rect -417 -185 -410 -180
rect -417 -187 -414 -185
rect -412 -187 -410 -185
rect -417 -189 -410 -187
rect -417 -194 -412 -189
rect -403 -191 -394 -174
rect -403 -193 -400 -191
rect -398 -192 -394 -191
rect -392 -176 -385 -174
rect -392 -178 -389 -176
rect -387 -178 -385 -176
rect -392 -183 -385 -178
rect -392 -185 -389 -183
rect -387 -185 -385 -183
rect -392 -187 -385 -185
rect -392 -192 -387 -187
rect -377 -191 -368 -174
rect -398 -193 -396 -192
rect -573 -205 -567 -203
rect -447 -201 -441 -194
rect -403 -195 -396 -193
rect -377 -193 -374 -191
rect -372 -192 -368 -191
rect -366 -176 -359 -174
rect -366 -178 -363 -176
rect -361 -178 -359 -176
rect -366 -183 -359 -178
rect -366 -185 -363 -183
rect -361 -185 -359 -183
rect -366 -187 -359 -185
rect -353 -182 -346 -180
rect -353 -184 -351 -182
rect -349 -184 -346 -182
rect -366 -192 -361 -187
rect -353 -189 -346 -184
rect -353 -191 -351 -189
rect -349 -191 -346 -189
rect -372 -193 -370 -192
rect -377 -195 -370 -193
rect -353 -193 -346 -191
rect -344 -181 -339 -180
rect -320 -181 -314 -176
rect -344 -193 -334 -181
rect -342 -194 -334 -193
rect -332 -183 -324 -181
rect -332 -185 -329 -183
rect -327 -185 -324 -183
rect -332 -190 -324 -185
rect -332 -192 -329 -190
rect -327 -192 -324 -190
rect -332 -194 -324 -192
rect -322 -190 -314 -181
rect -322 -192 -319 -190
rect -317 -192 -314 -190
rect -322 -194 -314 -192
rect -312 -178 -305 -176
rect -312 -180 -309 -178
rect -307 -180 -305 -178
rect -312 -185 -305 -180
rect -312 -187 -309 -185
rect -307 -187 -305 -185
rect -312 -189 -305 -187
rect -299 -182 -292 -180
rect -299 -184 -297 -182
rect -295 -184 -292 -182
rect -299 -189 -292 -184
rect -312 -194 -307 -189
rect -299 -191 -297 -189
rect -295 -191 -292 -189
rect -299 -193 -292 -191
rect -290 -181 -285 -180
rect -266 -181 -260 -176
rect -290 -193 -280 -181
rect -447 -203 -445 -201
rect -443 -203 -441 -201
rect -447 -205 -441 -203
rect -342 -201 -336 -194
rect -288 -194 -280 -193
rect -278 -183 -270 -181
rect -278 -185 -275 -183
rect -273 -185 -270 -183
rect -278 -190 -270 -185
rect -278 -192 -275 -190
rect -273 -192 -270 -190
rect -278 -194 -270 -192
rect -268 -190 -260 -181
rect -268 -192 -265 -190
rect -263 -192 -260 -190
rect -268 -194 -260 -192
rect -258 -178 -251 -176
rect -258 -180 -255 -178
rect -253 -180 -251 -178
rect -258 -185 -251 -180
rect -258 -187 -255 -185
rect -253 -187 -251 -185
rect -258 -189 -251 -187
rect -258 -194 -253 -189
rect -245 -191 -236 -174
rect -245 -193 -243 -191
rect -241 -193 -236 -191
rect -342 -203 -340 -201
rect -338 -203 -336 -201
rect -342 -205 -336 -203
rect -288 -201 -282 -194
rect -245 -198 -236 -193
rect -288 -203 -286 -201
rect -284 -203 -282 -201
rect -245 -200 -243 -198
rect -241 -200 -236 -198
rect -245 -202 -236 -200
rect -234 -202 -229 -174
rect -227 -182 -222 -174
rect -227 -184 -220 -182
rect -227 -186 -224 -184
rect -222 -186 -220 -184
rect -227 -191 -220 -186
rect -227 -193 -224 -191
rect -222 -193 -220 -191
rect -227 -195 -220 -193
rect -210 -191 -201 -174
rect -210 -193 -208 -191
rect -206 -193 -201 -191
rect -227 -202 -222 -195
rect -210 -198 -201 -193
rect -210 -200 -208 -198
rect -206 -200 -201 -198
rect -210 -202 -201 -200
rect -199 -202 -194 -174
rect -192 -182 -187 -174
rect -173 -182 -166 -180
rect -192 -184 -185 -182
rect -192 -186 -189 -184
rect -187 -186 -185 -184
rect -192 -191 -185 -186
rect -192 -193 -189 -191
rect -187 -193 -185 -191
rect -173 -184 -171 -182
rect -169 -184 -166 -182
rect -173 -189 -166 -184
rect -173 -191 -171 -189
rect -169 -191 -166 -189
rect -173 -193 -166 -191
rect -164 -181 -159 -180
rect -140 -181 -134 -176
rect -164 -193 -154 -181
rect -192 -195 -185 -193
rect -192 -202 -187 -195
rect -162 -194 -154 -193
rect -152 -183 -144 -181
rect -152 -185 -149 -183
rect -147 -185 -144 -183
rect -152 -190 -144 -185
rect -152 -192 -149 -190
rect -147 -192 -144 -190
rect -152 -194 -144 -192
rect -142 -190 -134 -181
rect -142 -192 -139 -190
rect -137 -192 -134 -190
rect -142 -194 -134 -192
rect -132 -178 -125 -176
rect -132 -180 -129 -178
rect -127 -180 -125 -178
rect -132 -185 -125 -180
rect -132 -187 -129 -185
rect -127 -187 -125 -185
rect -132 -189 -125 -187
rect -132 -194 -127 -189
rect -118 -191 -109 -174
rect -118 -193 -115 -191
rect -113 -192 -109 -191
rect -107 -176 -100 -174
rect -107 -178 -104 -176
rect -102 -178 -100 -176
rect -107 -183 -100 -178
rect -107 -185 -104 -183
rect -102 -185 -100 -183
rect -107 -187 -100 -185
rect -107 -192 -102 -187
rect -92 -191 -83 -174
rect -113 -193 -111 -192
rect -288 -205 -282 -203
rect -162 -201 -156 -194
rect -118 -195 -111 -193
rect -92 -193 -89 -191
rect -87 -192 -83 -191
rect -81 -176 -74 -174
rect -81 -178 -78 -176
rect -76 -178 -74 -176
rect -81 -183 -74 -178
rect -81 -185 -78 -183
rect -76 -185 -74 -183
rect -81 -187 -74 -185
rect -68 -182 -61 -180
rect -68 -184 -66 -182
rect -64 -184 -61 -182
rect -81 -192 -76 -187
rect -68 -189 -61 -184
rect -68 -191 -66 -189
rect -64 -191 -61 -189
rect -87 -193 -85 -192
rect -92 -195 -85 -193
rect -68 -193 -61 -191
rect -59 -181 -54 -180
rect -35 -181 -29 -176
rect -59 -193 -49 -181
rect -57 -194 -49 -193
rect -47 -183 -39 -181
rect -47 -185 -44 -183
rect -42 -185 -39 -183
rect -47 -190 -39 -185
rect -47 -192 -44 -190
rect -42 -192 -39 -190
rect -47 -194 -39 -192
rect -37 -190 -29 -181
rect -37 -192 -34 -190
rect -32 -192 -29 -190
rect -37 -194 -29 -192
rect -27 -178 -20 -176
rect -27 -180 -24 -178
rect -22 -180 -20 -178
rect -27 -185 -20 -180
rect -27 -187 -24 -185
rect -22 -187 -20 -185
rect -27 -189 -20 -187
rect -14 -182 -7 -180
rect -14 -184 -12 -182
rect -10 -184 -7 -182
rect -14 -189 -7 -184
rect -27 -194 -22 -189
rect -14 -191 -12 -189
rect -10 -191 -7 -189
rect -14 -193 -7 -191
rect -5 -181 0 -180
rect 19 -181 25 -176
rect -5 -193 5 -181
rect -162 -203 -160 -201
rect -158 -203 -156 -201
rect -162 -205 -156 -203
rect -57 -201 -51 -194
rect -3 -194 5 -193
rect 7 -183 15 -181
rect 7 -185 10 -183
rect 12 -185 15 -183
rect 7 -190 15 -185
rect 7 -192 10 -190
rect 12 -192 15 -190
rect 7 -194 15 -192
rect 17 -190 25 -181
rect 17 -192 20 -190
rect 22 -192 25 -190
rect 17 -194 25 -192
rect 27 -178 34 -176
rect 27 -180 30 -178
rect 32 -180 34 -178
rect 27 -185 34 -180
rect 27 -187 30 -185
rect 32 -187 34 -185
rect 27 -189 34 -187
rect 27 -194 32 -189
rect 40 -191 49 -174
rect 40 -193 42 -191
rect 44 -193 49 -191
rect -57 -203 -55 -201
rect -53 -203 -51 -201
rect -57 -205 -51 -203
rect -3 -201 3 -194
rect 40 -198 49 -193
rect -3 -203 -1 -201
rect 1 -203 3 -201
rect 40 -200 42 -198
rect 44 -200 49 -198
rect 40 -202 49 -200
rect 51 -202 56 -174
rect 58 -182 63 -174
rect 58 -184 65 -182
rect 58 -186 61 -184
rect 63 -186 65 -184
rect 58 -191 65 -186
rect 58 -193 61 -191
rect 63 -193 65 -191
rect 58 -195 65 -193
rect 75 -191 84 -174
rect 75 -193 77 -191
rect 79 -193 84 -191
rect 58 -202 63 -195
rect 75 -198 84 -193
rect 75 -200 77 -198
rect 79 -200 84 -198
rect 75 -202 84 -200
rect 86 -202 91 -174
rect 93 -182 98 -174
rect 112 -182 119 -180
rect 93 -184 100 -182
rect 93 -186 96 -184
rect 98 -186 100 -184
rect 93 -191 100 -186
rect 93 -193 96 -191
rect 98 -193 100 -191
rect 112 -184 114 -182
rect 116 -184 119 -182
rect 112 -189 119 -184
rect 112 -191 114 -189
rect 116 -191 119 -189
rect 112 -193 119 -191
rect 121 -181 126 -180
rect 145 -181 151 -176
rect 121 -193 131 -181
rect 93 -195 100 -193
rect 93 -202 98 -195
rect 123 -194 131 -193
rect 133 -183 141 -181
rect 133 -185 136 -183
rect 138 -185 141 -183
rect 133 -190 141 -185
rect 133 -192 136 -190
rect 138 -192 141 -190
rect 133 -194 141 -192
rect 143 -190 151 -181
rect 143 -192 146 -190
rect 148 -192 151 -190
rect 143 -194 151 -192
rect 153 -178 160 -176
rect 153 -180 156 -178
rect 158 -180 160 -178
rect 153 -185 160 -180
rect 153 -187 156 -185
rect 158 -187 160 -185
rect 153 -189 160 -187
rect 153 -194 158 -189
rect 167 -191 176 -174
rect 167 -193 170 -191
rect 172 -192 176 -191
rect 178 -176 185 -174
rect 178 -178 181 -176
rect 183 -178 185 -176
rect 178 -183 185 -178
rect 178 -185 181 -183
rect 183 -185 185 -183
rect 178 -187 185 -185
rect 178 -192 183 -187
rect 193 -191 202 -174
rect 172 -193 174 -192
rect -3 -205 3 -203
rect 123 -201 129 -194
rect 167 -195 174 -193
rect 193 -193 196 -191
rect 198 -192 202 -191
rect 204 -176 211 -174
rect 204 -178 207 -176
rect 209 -178 211 -176
rect 204 -183 211 -178
rect 204 -185 207 -183
rect 209 -185 211 -183
rect 204 -187 211 -185
rect 217 -182 224 -180
rect 217 -184 219 -182
rect 221 -184 224 -182
rect 204 -192 209 -187
rect 217 -189 224 -184
rect 217 -191 219 -189
rect 221 -191 224 -189
rect 198 -193 200 -192
rect 193 -195 200 -193
rect 217 -193 224 -191
rect 226 -181 231 -180
rect 250 -181 256 -176
rect 226 -193 236 -181
rect 228 -194 236 -193
rect 238 -183 246 -181
rect 238 -185 241 -183
rect 243 -185 246 -183
rect 238 -190 246 -185
rect 238 -192 241 -190
rect 243 -192 246 -190
rect 238 -194 246 -192
rect 248 -190 256 -181
rect 248 -192 251 -190
rect 253 -192 256 -190
rect 248 -194 256 -192
rect 258 -178 265 -176
rect 258 -180 261 -178
rect 263 -180 265 -178
rect 258 -185 265 -180
rect 258 -187 261 -185
rect 263 -187 265 -185
rect 258 -189 265 -187
rect 271 -182 278 -180
rect 271 -184 273 -182
rect 275 -184 278 -182
rect 271 -189 278 -184
rect 258 -194 263 -189
rect 271 -191 273 -189
rect 275 -191 278 -189
rect 271 -193 278 -191
rect 280 -181 285 -180
rect 304 -181 310 -176
rect 280 -193 290 -181
rect 123 -203 125 -201
rect 127 -203 129 -201
rect 123 -205 129 -203
rect 228 -201 234 -194
rect 282 -194 290 -193
rect 292 -183 300 -181
rect 292 -185 295 -183
rect 297 -185 300 -183
rect 292 -190 300 -185
rect 292 -192 295 -190
rect 297 -192 300 -190
rect 292 -194 300 -192
rect 302 -190 310 -181
rect 302 -192 305 -190
rect 307 -192 310 -190
rect 302 -194 310 -192
rect 312 -178 319 -176
rect 312 -180 315 -178
rect 317 -180 319 -178
rect 312 -185 319 -180
rect 312 -187 315 -185
rect 317 -187 319 -185
rect 312 -189 319 -187
rect 312 -194 317 -189
rect 325 -191 334 -174
rect 325 -193 327 -191
rect 329 -193 334 -191
rect 228 -203 230 -201
rect 232 -203 234 -201
rect 228 -205 234 -203
rect 282 -201 288 -194
rect 325 -198 334 -193
rect 282 -203 284 -201
rect 286 -203 288 -201
rect 325 -200 327 -198
rect 329 -200 334 -198
rect 325 -202 334 -200
rect 336 -202 341 -174
rect 343 -182 348 -174
rect 343 -184 350 -182
rect 343 -186 346 -184
rect 348 -186 350 -184
rect 343 -191 350 -186
rect 343 -193 346 -191
rect 348 -193 350 -191
rect 343 -195 350 -193
rect 360 -191 369 -174
rect 360 -193 362 -191
rect 364 -193 369 -191
rect 343 -202 348 -195
rect 360 -198 369 -193
rect 360 -200 362 -198
rect 364 -200 369 -198
rect 360 -202 369 -200
rect 371 -202 376 -174
rect 378 -182 383 -174
rect 397 -182 404 -180
rect 378 -184 385 -182
rect 378 -186 381 -184
rect 383 -186 385 -184
rect 378 -191 385 -186
rect 378 -193 381 -191
rect 383 -193 385 -191
rect 397 -184 399 -182
rect 401 -184 404 -182
rect 397 -189 404 -184
rect 397 -191 399 -189
rect 401 -191 404 -189
rect 397 -193 404 -191
rect 406 -181 411 -180
rect 430 -181 436 -176
rect 406 -193 416 -181
rect 378 -195 385 -193
rect 378 -202 383 -195
rect 408 -194 416 -193
rect 418 -183 426 -181
rect 418 -185 421 -183
rect 423 -185 426 -183
rect 418 -190 426 -185
rect 418 -192 421 -190
rect 423 -192 426 -190
rect 418 -194 426 -192
rect 428 -190 436 -181
rect 428 -192 431 -190
rect 433 -192 436 -190
rect 428 -194 436 -192
rect 438 -178 445 -176
rect 438 -180 441 -178
rect 443 -180 445 -178
rect 438 -185 445 -180
rect 524 -182 529 -174
rect 438 -187 441 -185
rect 443 -187 445 -185
rect 438 -189 445 -187
rect 438 -194 443 -189
rect 282 -205 288 -203
rect 408 -201 414 -194
rect 458 -196 465 -182
rect 458 -198 460 -196
rect 462 -198 465 -196
rect 458 -200 465 -198
rect 467 -200 472 -182
rect 474 -200 479 -182
rect 481 -200 486 -182
rect 488 -191 496 -182
rect 488 -193 491 -191
rect 493 -193 496 -191
rect 488 -200 496 -193
rect 498 -200 503 -182
rect 505 -200 510 -182
rect 512 -200 517 -182
rect 519 -192 529 -182
rect 531 -176 538 -174
rect 531 -178 534 -176
rect 536 -178 538 -176
rect 531 -183 538 -178
rect 616 -182 621 -174
rect 531 -185 534 -183
rect 536 -185 538 -183
rect 531 -187 538 -185
rect 531 -192 536 -187
rect 519 -198 527 -192
rect 550 -196 557 -182
rect 519 -200 523 -198
rect 525 -200 527 -198
rect 550 -198 552 -196
rect 554 -198 557 -196
rect 408 -203 410 -201
rect 412 -203 414 -201
rect 408 -205 414 -203
rect 521 -202 527 -200
rect 550 -200 557 -198
rect 559 -200 564 -182
rect 566 -200 571 -182
rect 573 -200 578 -182
rect 580 -191 588 -182
rect 580 -193 583 -191
rect 585 -193 588 -191
rect 580 -200 588 -193
rect 590 -200 595 -182
rect 597 -200 602 -182
rect 604 -200 609 -182
rect 611 -192 621 -182
rect 623 -176 630 -174
rect 623 -178 626 -176
rect 628 -178 630 -176
rect 623 -183 630 -178
rect 623 -185 626 -183
rect 628 -185 630 -183
rect 623 -187 630 -185
rect 623 -192 628 -187
rect 611 -198 619 -192
rect 611 -200 615 -198
rect 617 -200 619 -198
rect 613 -202 619 -200
rect -627 -213 -621 -211
rect -627 -215 -625 -213
rect -623 -215 -621 -213
rect -688 -223 -681 -221
rect -688 -225 -685 -223
rect -683 -224 -681 -223
rect -662 -223 -655 -221
rect -683 -225 -679 -224
rect -688 -242 -679 -225
rect -677 -229 -672 -224
rect -662 -225 -659 -223
rect -657 -224 -655 -223
rect -627 -222 -621 -215
rect -573 -213 -567 -211
rect -573 -215 -571 -213
rect -569 -215 -567 -213
rect -627 -223 -619 -222
rect -657 -225 -653 -224
rect -677 -231 -670 -229
rect -677 -233 -674 -231
rect -672 -233 -670 -231
rect -677 -238 -670 -233
rect -677 -240 -674 -238
rect -672 -240 -670 -238
rect -677 -242 -670 -240
rect -662 -242 -653 -225
rect -651 -229 -646 -224
rect -638 -225 -631 -223
rect -638 -227 -636 -225
rect -634 -227 -631 -225
rect -651 -231 -644 -229
rect -651 -233 -648 -231
rect -646 -233 -644 -231
rect -651 -238 -644 -233
rect -638 -232 -631 -227
rect -638 -234 -636 -232
rect -634 -234 -631 -232
rect -638 -236 -631 -234
rect -629 -235 -619 -223
rect -617 -224 -609 -222
rect -617 -226 -614 -224
rect -612 -226 -609 -224
rect -617 -231 -609 -226
rect -617 -233 -614 -231
rect -612 -233 -609 -231
rect -617 -235 -609 -233
rect -607 -224 -599 -222
rect -607 -226 -604 -224
rect -602 -226 -599 -224
rect -607 -235 -599 -226
rect -629 -236 -624 -235
rect -651 -240 -648 -238
rect -646 -240 -644 -238
rect -651 -242 -644 -240
rect -605 -240 -599 -235
rect -597 -227 -592 -222
rect -573 -222 -567 -215
rect -530 -216 -521 -214
rect -530 -218 -528 -216
rect -526 -218 -521 -216
rect -573 -223 -565 -222
rect -584 -225 -577 -223
rect -584 -227 -582 -225
rect -580 -227 -577 -225
rect -597 -229 -590 -227
rect -597 -231 -594 -229
rect -592 -231 -590 -229
rect -597 -236 -590 -231
rect -584 -232 -577 -227
rect -584 -234 -582 -232
rect -580 -234 -577 -232
rect -584 -236 -577 -234
rect -575 -235 -565 -223
rect -563 -224 -555 -222
rect -563 -226 -560 -224
rect -558 -226 -555 -224
rect -563 -231 -555 -226
rect -563 -233 -560 -231
rect -558 -233 -555 -231
rect -563 -235 -555 -233
rect -553 -224 -545 -222
rect -553 -226 -550 -224
rect -548 -226 -545 -224
rect -553 -235 -545 -226
rect -575 -236 -570 -235
rect -597 -238 -594 -236
rect -592 -238 -590 -236
rect -597 -240 -590 -238
rect -551 -240 -545 -235
rect -543 -227 -538 -222
rect -530 -223 -521 -218
rect -530 -225 -528 -223
rect -526 -225 -521 -223
rect -543 -229 -536 -227
rect -543 -231 -540 -229
rect -538 -231 -536 -229
rect -543 -236 -536 -231
rect -543 -238 -540 -236
rect -538 -238 -536 -236
rect -543 -240 -536 -238
rect -530 -242 -521 -225
rect -519 -242 -514 -214
rect -512 -221 -507 -214
rect -495 -216 -486 -214
rect -495 -218 -493 -216
rect -491 -218 -486 -216
rect -512 -223 -505 -221
rect -512 -225 -509 -223
rect -507 -225 -505 -223
rect -512 -230 -505 -225
rect -512 -232 -509 -230
rect -507 -232 -505 -230
rect -512 -234 -505 -232
rect -495 -223 -486 -218
rect -495 -225 -493 -223
rect -491 -225 -486 -223
rect -512 -242 -507 -234
rect -495 -242 -486 -225
rect -484 -242 -479 -214
rect -477 -221 -472 -214
rect -447 -213 -441 -211
rect -447 -215 -445 -213
rect -443 -215 -441 -213
rect -477 -223 -470 -221
rect -447 -222 -441 -215
rect -342 -213 -336 -211
rect -342 -215 -340 -213
rect -338 -215 -336 -213
rect -447 -223 -439 -222
rect -477 -225 -474 -223
rect -472 -225 -470 -223
rect -477 -230 -470 -225
rect -477 -232 -474 -230
rect -472 -232 -470 -230
rect -477 -234 -470 -232
rect -458 -225 -451 -223
rect -458 -227 -456 -225
rect -454 -227 -451 -225
rect -458 -232 -451 -227
rect -458 -234 -456 -232
rect -454 -234 -451 -232
rect -477 -242 -472 -234
rect -458 -236 -451 -234
rect -449 -235 -439 -223
rect -437 -224 -429 -222
rect -437 -226 -434 -224
rect -432 -226 -429 -224
rect -437 -231 -429 -226
rect -437 -233 -434 -231
rect -432 -233 -429 -231
rect -437 -235 -429 -233
rect -427 -224 -419 -222
rect -427 -226 -424 -224
rect -422 -226 -419 -224
rect -427 -235 -419 -226
rect -449 -236 -444 -235
rect -425 -240 -419 -235
rect -417 -227 -412 -222
rect -403 -223 -396 -221
rect -403 -225 -400 -223
rect -398 -224 -396 -223
rect -377 -223 -370 -221
rect -398 -225 -394 -224
rect -417 -229 -410 -227
rect -417 -231 -414 -229
rect -412 -231 -410 -229
rect -417 -236 -410 -231
rect -417 -238 -414 -236
rect -412 -238 -410 -236
rect -417 -240 -410 -238
rect -403 -242 -394 -225
rect -392 -229 -387 -224
rect -377 -225 -374 -223
rect -372 -224 -370 -223
rect -342 -222 -336 -215
rect -288 -213 -282 -211
rect -288 -215 -286 -213
rect -284 -215 -282 -213
rect -342 -223 -334 -222
rect -372 -225 -368 -224
rect -392 -231 -385 -229
rect -392 -233 -389 -231
rect -387 -233 -385 -231
rect -392 -238 -385 -233
rect -392 -240 -389 -238
rect -387 -240 -385 -238
rect -392 -242 -385 -240
rect -377 -242 -368 -225
rect -366 -229 -361 -224
rect -353 -225 -346 -223
rect -353 -227 -351 -225
rect -349 -227 -346 -225
rect -366 -231 -359 -229
rect -366 -233 -363 -231
rect -361 -233 -359 -231
rect -366 -238 -359 -233
rect -353 -232 -346 -227
rect -353 -234 -351 -232
rect -349 -234 -346 -232
rect -353 -236 -346 -234
rect -344 -235 -334 -223
rect -332 -224 -324 -222
rect -332 -226 -329 -224
rect -327 -226 -324 -224
rect -332 -231 -324 -226
rect -332 -233 -329 -231
rect -327 -233 -324 -231
rect -332 -235 -324 -233
rect -322 -224 -314 -222
rect -322 -226 -319 -224
rect -317 -226 -314 -224
rect -322 -235 -314 -226
rect -344 -236 -339 -235
rect -366 -240 -363 -238
rect -361 -240 -359 -238
rect -366 -242 -359 -240
rect -320 -240 -314 -235
rect -312 -227 -307 -222
rect -288 -222 -282 -215
rect -245 -216 -236 -214
rect -245 -218 -243 -216
rect -241 -218 -236 -216
rect -288 -223 -280 -222
rect -299 -225 -292 -223
rect -299 -227 -297 -225
rect -295 -227 -292 -225
rect -312 -229 -305 -227
rect -312 -231 -309 -229
rect -307 -231 -305 -229
rect -312 -236 -305 -231
rect -299 -232 -292 -227
rect -299 -234 -297 -232
rect -295 -234 -292 -232
rect -299 -236 -292 -234
rect -290 -235 -280 -223
rect -278 -224 -270 -222
rect -278 -226 -275 -224
rect -273 -226 -270 -224
rect -278 -231 -270 -226
rect -278 -233 -275 -231
rect -273 -233 -270 -231
rect -278 -235 -270 -233
rect -268 -224 -260 -222
rect -268 -226 -265 -224
rect -263 -226 -260 -224
rect -268 -235 -260 -226
rect -290 -236 -285 -235
rect -312 -238 -309 -236
rect -307 -238 -305 -236
rect -312 -240 -305 -238
rect -266 -240 -260 -235
rect -258 -227 -253 -222
rect -245 -223 -236 -218
rect -245 -225 -243 -223
rect -241 -225 -236 -223
rect -258 -229 -251 -227
rect -258 -231 -255 -229
rect -253 -231 -251 -229
rect -258 -236 -251 -231
rect -258 -238 -255 -236
rect -253 -238 -251 -236
rect -258 -240 -251 -238
rect -245 -242 -236 -225
rect -234 -242 -229 -214
rect -227 -221 -222 -214
rect -210 -216 -201 -214
rect -210 -218 -208 -216
rect -206 -218 -201 -216
rect -227 -223 -220 -221
rect -227 -225 -224 -223
rect -222 -225 -220 -223
rect -227 -230 -220 -225
rect -227 -232 -224 -230
rect -222 -232 -220 -230
rect -227 -234 -220 -232
rect -210 -223 -201 -218
rect -210 -225 -208 -223
rect -206 -225 -201 -223
rect -227 -242 -222 -234
rect -210 -242 -201 -225
rect -199 -242 -194 -214
rect -192 -221 -187 -214
rect -162 -213 -156 -211
rect -162 -215 -160 -213
rect -158 -215 -156 -213
rect -192 -223 -185 -221
rect -162 -222 -156 -215
rect -57 -213 -51 -211
rect -57 -215 -55 -213
rect -53 -215 -51 -213
rect -162 -223 -154 -222
rect -192 -225 -189 -223
rect -187 -225 -185 -223
rect -192 -230 -185 -225
rect -192 -232 -189 -230
rect -187 -232 -185 -230
rect -192 -234 -185 -232
rect -173 -225 -166 -223
rect -173 -227 -171 -225
rect -169 -227 -166 -225
rect -173 -232 -166 -227
rect -173 -234 -171 -232
rect -169 -234 -166 -232
rect -192 -242 -187 -234
rect -173 -236 -166 -234
rect -164 -235 -154 -223
rect -152 -224 -144 -222
rect -152 -226 -149 -224
rect -147 -226 -144 -224
rect -152 -231 -144 -226
rect -152 -233 -149 -231
rect -147 -233 -144 -231
rect -152 -235 -144 -233
rect -142 -224 -134 -222
rect -142 -226 -139 -224
rect -137 -226 -134 -224
rect -142 -235 -134 -226
rect -164 -236 -159 -235
rect -140 -240 -134 -235
rect -132 -227 -127 -222
rect -118 -223 -111 -221
rect -118 -225 -115 -223
rect -113 -224 -111 -223
rect -92 -223 -85 -221
rect -113 -225 -109 -224
rect -132 -229 -125 -227
rect -132 -231 -129 -229
rect -127 -231 -125 -229
rect -132 -236 -125 -231
rect -132 -238 -129 -236
rect -127 -238 -125 -236
rect -132 -240 -125 -238
rect -118 -242 -109 -225
rect -107 -229 -102 -224
rect -92 -225 -89 -223
rect -87 -224 -85 -223
rect -57 -222 -51 -215
rect -3 -213 3 -211
rect -3 -215 -1 -213
rect 1 -215 3 -213
rect -57 -223 -49 -222
rect -87 -225 -83 -224
rect -107 -231 -100 -229
rect -107 -233 -104 -231
rect -102 -233 -100 -231
rect -107 -238 -100 -233
rect -107 -240 -104 -238
rect -102 -240 -100 -238
rect -107 -242 -100 -240
rect -92 -242 -83 -225
rect -81 -229 -76 -224
rect -68 -225 -61 -223
rect -68 -227 -66 -225
rect -64 -227 -61 -225
rect -81 -231 -74 -229
rect -81 -233 -78 -231
rect -76 -233 -74 -231
rect -81 -238 -74 -233
rect -68 -232 -61 -227
rect -68 -234 -66 -232
rect -64 -234 -61 -232
rect -68 -236 -61 -234
rect -59 -235 -49 -223
rect -47 -224 -39 -222
rect -47 -226 -44 -224
rect -42 -226 -39 -224
rect -47 -231 -39 -226
rect -47 -233 -44 -231
rect -42 -233 -39 -231
rect -47 -235 -39 -233
rect -37 -224 -29 -222
rect -37 -226 -34 -224
rect -32 -226 -29 -224
rect -37 -235 -29 -226
rect -59 -236 -54 -235
rect -81 -240 -78 -238
rect -76 -240 -74 -238
rect -81 -242 -74 -240
rect -35 -240 -29 -235
rect -27 -227 -22 -222
rect -3 -222 3 -215
rect 40 -216 49 -214
rect 40 -218 42 -216
rect 44 -218 49 -216
rect -3 -223 5 -222
rect -14 -225 -7 -223
rect -14 -227 -12 -225
rect -10 -227 -7 -225
rect -27 -229 -20 -227
rect -27 -231 -24 -229
rect -22 -231 -20 -229
rect -27 -236 -20 -231
rect -14 -232 -7 -227
rect -14 -234 -12 -232
rect -10 -234 -7 -232
rect -14 -236 -7 -234
rect -5 -235 5 -223
rect 7 -224 15 -222
rect 7 -226 10 -224
rect 12 -226 15 -224
rect 7 -231 15 -226
rect 7 -233 10 -231
rect 12 -233 15 -231
rect 7 -235 15 -233
rect 17 -224 25 -222
rect 17 -226 20 -224
rect 22 -226 25 -224
rect 17 -235 25 -226
rect -5 -236 0 -235
rect -27 -238 -24 -236
rect -22 -238 -20 -236
rect -27 -240 -20 -238
rect 19 -240 25 -235
rect 27 -227 32 -222
rect 40 -223 49 -218
rect 40 -225 42 -223
rect 44 -225 49 -223
rect 27 -229 34 -227
rect 27 -231 30 -229
rect 32 -231 34 -229
rect 27 -236 34 -231
rect 27 -238 30 -236
rect 32 -238 34 -236
rect 27 -240 34 -238
rect 40 -242 49 -225
rect 51 -242 56 -214
rect 58 -221 63 -214
rect 75 -216 84 -214
rect 75 -218 77 -216
rect 79 -218 84 -216
rect 58 -223 65 -221
rect 58 -225 61 -223
rect 63 -225 65 -223
rect 58 -230 65 -225
rect 58 -232 61 -230
rect 63 -232 65 -230
rect 58 -234 65 -232
rect 75 -223 84 -218
rect 75 -225 77 -223
rect 79 -225 84 -223
rect 58 -242 63 -234
rect 75 -242 84 -225
rect 86 -242 91 -214
rect 93 -221 98 -214
rect 123 -213 129 -211
rect 123 -215 125 -213
rect 127 -215 129 -213
rect 93 -223 100 -221
rect 123 -222 129 -215
rect 228 -213 234 -211
rect 228 -215 230 -213
rect 232 -215 234 -213
rect 123 -223 131 -222
rect 93 -225 96 -223
rect 98 -225 100 -223
rect 93 -230 100 -225
rect 93 -232 96 -230
rect 98 -232 100 -230
rect 93 -234 100 -232
rect 112 -225 119 -223
rect 112 -227 114 -225
rect 116 -227 119 -225
rect 112 -232 119 -227
rect 112 -234 114 -232
rect 116 -234 119 -232
rect 93 -242 98 -234
rect 112 -236 119 -234
rect 121 -235 131 -223
rect 133 -224 141 -222
rect 133 -226 136 -224
rect 138 -226 141 -224
rect 133 -231 141 -226
rect 133 -233 136 -231
rect 138 -233 141 -231
rect 133 -235 141 -233
rect 143 -224 151 -222
rect 143 -226 146 -224
rect 148 -226 151 -224
rect 143 -235 151 -226
rect 121 -236 126 -235
rect 145 -240 151 -235
rect 153 -227 158 -222
rect 167 -223 174 -221
rect 167 -225 170 -223
rect 172 -224 174 -223
rect 193 -223 200 -221
rect 172 -225 176 -224
rect 153 -229 160 -227
rect 153 -231 156 -229
rect 158 -231 160 -229
rect 153 -236 160 -231
rect 153 -238 156 -236
rect 158 -238 160 -236
rect 153 -240 160 -238
rect 167 -242 176 -225
rect 178 -229 183 -224
rect 193 -225 196 -223
rect 198 -224 200 -223
rect 228 -222 234 -215
rect 282 -213 288 -211
rect 282 -215 284 -213
rect 286 -215 288 -213
rect 228 -223 236 -222
rect 198 -225 202 -224
rect 178 -231 185 -229
rect 178 -233 181 -231
rect 183 -233 185 -231
rect 178 -238 185 -233
rect 178 -240 181 -238
rect 183 -240 185 -238
rect 178 -242 185 -240
rect 193 -242 202 -225
rect 204 -229 209 -224
rect 217 -225 224 -223
rect 217 -227 219 -225
rect 221 -227 224 -225
rect 204 -231 211 -229
rect 204 -233 207 -231
rect 209 -233 211 -231
rect 204 -238 211 -233
rect 217 -232 224 -227
rect 217 -234 219 -232
rect 221 -234 224 -232
rect 217 -236 224 -234
rect 226 -235 236 -223
rect 238 -224 246 -222
rect 238 -226 241 -224
rect 243 -226 246 -224
rect 238 -231 246 -226
rect 238 -233 241 -231
rect 243 -233 246 -231
rect 238 -235 246 -233
rect 248 -224 256 -222
rect 248 -226 251 -224
rect 253 -226 256 -224
rect 248 -235 256 -226
rect 226 -236 231 -235
rect 204 -240 207 -238
rect 209 -240 211 -238
rect 204 -242 211 -240
rect 250 -240 256 -235
rect 258 -227 263 -222
rect 282 -222 288 -215
rect 325 -216 334 -214
rect 325 -218 327 -216
rect 329 -218 334 -216
rect 282 -223 290 -222
rect 271 -225 278 -223
rect 271 -227 273 -225
rect 275 -227 278 -225
rect 258 -229 265 -227
rect 258 -231 261 -229
rect 263 -231 265 -229
rect 258 -236 265 -231
rect 271 -232 278 -227
rect 271 -234 273 -232
rect 275 -234 278 -232
rect 271 -236 278 -234
rect 280 -235 290 -223
rect 292 -224 300 -222
rect 292 -226 295 -224
rect 297 -226 300 -224
rect 292 -231 300 -226
rect 292 -233 295 -231
rect 297 -233 300 -231
rect 292 -235 300 -233
rect 302 -224 310 -222
rect 302 -226 305 -224
rect 307 -226 310 -224
rect 302 -235 310 -226
rect 280 -236 285 -235
rect 258 -238 261 -236
rect 263 -238 265 -236
rect 258 -240 265 -238
rect 304 -240 310 -235
rect 312 -227 317 -222
rect 325 -223 334 -218
rect 325 -225 327 -223
rect 329 -225 334 -223
rect 312 -229 319 -227
rect 312 -231 315 -229
rect 317 -231 319 -229
rect 312 -236 319 -231
rect 312 -238 315 -236
rect 317 -238 319 -236
rect 312 -240 319 -238
rect 325 -242 334 -225
rect 336 -242 341 -214
rect 343 -221 348 -214
rect 360 -216 369 -214
rect 360 -218 362 -216
rect 364 -218 369 -216
rect 343 -223 350 -221
rect 343 -225 346 -223
rect 348 -225 350 -223
rect 343 -230 350 -225
rect 343 -232 346 -230
rect 348 -232 350 -230
rect 343 -234 350 -232
rect 360 -223 369 -218
rect 360 -225 362 -223
rect 364 -225 369 -223
rect 343 -242 348 -234
rect 360 -242 369 -225
rect 371 -242 376 -214
rect 378 -221 383 -214
rect 408 -213 414 -211
rect 408 -215 410 -213
rect 412 -215 414 -213
rect 378 -223 385 -221
rect 408 -222 414 -215
rect 521 -216 527 -214
rect 458 -218 465 -216
rect 458 -220 460 -218
rect 462 -220 465 -218
rect 408 -223 416 -222
rect 378 -225 381 -223
rect 383 -225 385 -223
rect 378 -230 385 -225
rect 378 -232 381 -230
rect 383 -232 385 -230
rect 378 -234 385 -232
rect 397 -225 404 -223
rect 397 -227 399 -225
rect 401 -227 404 -225
rect 397 -232 404 -227
rect 397 -234 399 -232
rect 401 -234 404 -232
rect 378 -242 383 -234
rect 397 -236 404 -234
rect 406 -235 416 -223
rect 418 -224 426 -222
rect 418 -226 421 -224
rect 423 -226 426 -224
rect 418 -231 426 -226
rect 418 -233 421 -231
rect 423 -233 426 -231
rect 418 -235 426 -233
rect 428 -224 436 -222
rect 428 -226 431 -224
rect 433 -226 436 -224
rect 428 -235 436 -226
rect 406 -236 411 -235
rect 430 -240 436 -235
rect 438 -227 443 -222
rect 438 -229 445 -227
rect 438 -231 441 -229
rect 443 -231 445 -229
rect 438 -236 445 -231
rect 458 -234 465 -220
rect 467 -234 472 -216
rect 474 -234 479 -216
rect 481 -234 486 -216
rect 488 -223 496 -216
rect 488 -225 491 -223
rect 493 -225 496 -223
rect 488 -234 496 -225
rect 498 -234 503 -216
rect 505 -234 510 -216
rect 512 -234 517 -216
rect 519 -218 523 -216
rect 525 -218 527 -216
rect 613 -216 619 -214
rect 519 -224 527 -218
rect 550 -218 557 -216
rect 550 -220 552 -218
rect 554 -220 557 -218
rect 519 -234 529 -224
rect 438 -238 441 -236
rect 443 -238 445 -236
rect 438 -240 445 -238
rect 524 -242 529 -234
rect 531 -229 536 -224
rect 531 -231 538 -229
rect 531 -233 534 -231
rect 536 -233 538 -231
rect 531 -238 538 -233
rect 550 -234 557 -220
rect 559 -234 564 -216
rect 566 -234 571 -216
rect 573 -234 578 -216
rect 580 -223 588 -216
rect 580 -225 583 -223
rect 585 -225 588 -223
rect 580 -234 588 -225
rect 590 -234 595 -216
rect 597 -234 602 -216
rect 604 -234 609 -216
rect 611 -218 615 -216
rect 617 -218 619 -216
rect 611 -224 619 -218
rect 611 -234 621 -224
rect 531 -240 534 -238
rect 536 -240 538 -238
rect 531 -242 538 -240
rect 616 -242 621 -234
rect 623 -229 628 -224
rect 623 -231 630 -229
rect 623 -233 626 -231
rect 628 -233 630 -231
rect 623 -238 630 -233
rect 623 -240 626 -238
rect 628 -240 630 -238
rect 623 -242 630 -240
<< alu1 >>
rect 178 318 676 319
rect 178 316 179 318
rect 181 316 673 318
rect 675 316 676 318
rect 178 315 676 316
rect 149 310 668 311
rect 149 308 150 310
rect 152 308 665 310
rect 667 308 668 310
rect 149 307 668 308
rect -104 302 153 303
rect -104 300 -103 302
rect -101 300 150 302
rect 152 300 153 302
rect -104 299 153 300
rect 157 302 660 303
rect 157 300 158 302
rect 160 300 657 302
rect 659 300 660 302
rect 157 299 660 300
rect -715 294 -685 295
rect -715 292 -714 294
rect -712 292 -688 294
rect -686 292 -685 294
rect -715 291 -685 292
rect -414 294 -123 295
rect -414 292 -413 294
rect -411 292 -126 294
rect -124 292 -123 294
rect -414 291 -123 292
rect -119 294 652 295
rect -119 292 -118 294
rect -116 292 649 294
rect 651 292 652 294
rect -119 291 652 292
rect -707 286 -400 287
rect -707 284 -706 286
rect -704 284 -403 286
rect -401 284 -400 286
rect -707 283 -400 284
rect -127 286 161 287
rect -127 284 -126 286
rect -124 284 158 286
rect 160 284 161 286
rect -127 283 161 284
rect 166 286 644 287
rect 166 284 167 286
rect 169 284 641 286
rect 643 284 644 286
rect 166 283 644 284
rect -664 278 195 279
rect -664 276 -663 278
rect -661 276 -378 278
rect -376 276 -93 278
rect -91 276 192 278
rect 194 276 195 278
rect -664 275 195 276
rect 441 278 684 279
rect 441 276 442 278
rect 444 276 681 278
rect 683 276 684 278
rect 441 275 684 276
rect -618 270 518 271
rect -618 268 -617 270
rect -615 268 -332 270
rect -330 268 -47 270
rect -45 268 238 270
rect 240 268 515 270
rect 517 268 518 270
rect -618 267 518 268
rect -618 262 -434 263
rect -618 260 -617 262
rect -615 260 -563 262
rect -561 260 -437 262
rect -435 260 -434 262
rect -618 259 -434 260
rect -333 262 -149 263
rect -333 260 -332 262
rect -330 260 -278 262
rect -276 260 -152 262
rect -150 260 -149 262
rect -333 259 -149 260
rect -48 262 136 263
rect -48 260 -47 262
rect -45 260 7 262
rect 9 260 133 262
rect 135 260 136 262
rect -48 259 136 260
rect 237 262 421 263
rect 237 260 238 262
rect 240 260 292 262
rect 294 260 418 262
rect 420 260 421 262
rect 237 259 421 260
rect 454 262 636 263
rect 454 260 455 262
rect 457 260 633 262
rect 635 260 636 262
rect 454 259 636 260
rect -664 254 -443 255
rect -664 252 -663 254
rect -661 252 -446 254
rect -444 252 -443 254
rect -664 251 -443 252
rect -379 254 -158 255
rect -379 252 -378 254
rect -376 252 -161 254
rect -159 252 -158 254
rect -379 251 -158 252
rect -94 254 127 255
rect -94 252 -93 254
rect -91 252 124 254
rect 126 252 127 254
rect -94 251 127 252
rect 191 254 412 255
rect 191 252 192 254
rect 194 252 409 254
rect 411 252 412 254
rect 191 251 412 252
rect 454 254 458 255
rect 454 252 455 254
rect 457 252 458 254
rect 454 251 458 252
rect 514 254 518 255
rect 514 252 515 254
rect 517 252 518 254
rect 514 251 518 252
rect -594 246 -479 247
rect -594 244 -593 246
rect -591 244 -482 246
rect -480 244 -479 246
rect -594 243 -479 244
rect -309 246 -194 247
rect -309 244 -308 246
rect -306 244 -197 246
rect -195 244 -194 246
rect -309 243 -194 244
rect -24 246 91 247
rect -24 244 -23 246
rect -21 244 88 246
rect 90 244 91 246
rect -24 243 91 244
rect 261 246 376 247
rect 261 244 262 246
rect 264 244 373 246
rect 375 244 376 246
rect 261 243 376 244
rect 478 246 612 247
rect 478 244 479 246
rect 481 244 539 246
rect 541 244 609 246
rect 611 244 612 246
rect 478 243 612 244
rect 156 242 182 243
rect 156 240 157 242
rect 159 240 179 242
rect 181 240 182 242
rect 156 239 182 240
rect -699 238 -660 239
rect -699 236 -698 238
rect -696 236 -663 238
rect -661 236 -660 238
rect -699 235 -660 236
rect -648 238 -569 239
rect -648 236 -647 238
rect -645 236 -626 238
rect -624 236 -572 238
rect -570 236 -569 238
rect -648 235 -569 236
rect -363 238 -284 239
rect -363 236 -362 238
rect -360 236 -341 238
rect -339 236 -287 238
rect -285 236 -284 238
rect -363 235 -284 236
rect -129 238 -100 239
rect -129 236 -128 238
rect -126 236 -103 238
rect -101 236 -100 238
rect -129 235 -100 236
rect -78 238 1 239
rect -78 236 -77 238
rect -75 236 -56 238
rect -54 236 -2 238
rect 0 236 1 238
rect -78 235 1 236
rect 207 238 286 239
rect 207 236 208 238
rect 210 236 229 238
rect 231 236 283 238
rect 285 236 286 238
rect 207 235 286 236
rect 550 238 628 239
rect 550 236 551 238
rect 553 236 581 238
rect 583 236 625 238
rect 627 236 628 238
rect 550 235 628 236
rect -689 230 -577 231
rect -689 228 -688 230
rect -686 228 -580 230
rect -578 228 -577 230
rect -689 227 -577 228
rect -514 230 -451 231
rect -514 228 -513 230
rect -511 228 -470 230
rect -468 228 -454 230
rect -452 228 -451 230
rect -514 227 -451 228
rect -404 230 -292 231
rect -404 228 -403 230
rect -401 228 -295 230
rect -293 228 -292 230
rect -404 227 -292 228
rect -229 230 -166 231
rect -229 228 -228 230
rect -226 228 -185 230
rect -183 228 -169 230
rect -167 228 -166 230
rect -229 227 -166 228
rect -119 230 -7 231
rect -119 228 -118 230
rect -116 228 -10 230
rect -8 228 -7 230
rect -119 227 -7 228
rect 56 230 119 231
rect 56 228 57 230
rect 59 228 100 230
rect 102 228 116 230
rect 118 228 119 230
rect 56 227 119 228
rect 166 230 278 231
rect 166 228 167 230
rect 169 228 275 230
rect 277 228 278 230
rect 166 227 278 228
rect 341 230 404 231
rect 341 228 342 230
rect 344 228 385 230
rect 387 228 401 230
rect 403 228 404 230
rect 341 227 404 228
rect 488 230 620 231
rect 488 228 489 230
rect 491 228 597 230
rect 599 228 617 230
rect 619 228 620 230
rect 488 227 620 228
rect -674 222 -631 223
rect -674 220 -673 222
rect -671 220 -634 222
rect -632 220 -631 222
rect -674 219 -631 220
rect -540 222 -526 223
rect -540 220 -539 222
rect -537 220 -529 222
rect -527 220 -526 222
rect -540 219 -526 220
rect -506 222 -491 223
rect -506 220 -505 222
rect -503 220 -494 222
rect -492 220 -491 222
rect -506 219 -491 220
rect -483 222 -479 223
rect -483 220 -482 222
rect -480 220 -479 222
rect -483 219 -479 220
rect -389 222 -346 223
rect -389 220 -388 222
rect -386 220 -349 222
rect -347 220 -346 222
rect -389 219 -346 220
rect -255 222 -241 223
rect -255 220 -254 222
rect -252 220 -244 222
rect -242 220 -241 222
rect -255 219 -241 220
rect -221 222 -206 223
rect -221 220 -220 222
rect -218 220 -209 222
rect -207 220 -206 222
rect -221 219 -206 220
rect -198 222 -194 223
rect -198 220 -197 222
rect -195 220 -194 222
rect -198 219 -194 220
rect -104 222 -61 223
rect -104 220 -103 222
rect -101 220 -64 222
rect -62 220 -61 222
rect -104 219 -61 220
rect 30 222 44 223
rect 30 220 31 222
rect 33 220 41 222
rect 43 220 44 222
rect 30 219 44 220
rect 64 222 79 223
rect 64 220 65 222
rect 67 220 76 222
rect 78 220 79 222
rect 64 219 79 220
rect 87 222 91 223
rect 87 220 88 222
rect 90 220 91 222
rect 87 219 91 220
rect 181 222 224 223
rect 181 220 182 222
rect 184 220 221 222
rect 223 220 224 222
rect 181 219 224 220
rect 315 222 329 223
rect 315 220 316 222
rect 318 220 326 222
rect 328 220 329 222
rect 315 219 329 220
rect 349 222 364 223
rect 349 220 350 222
rect 352 220 361 222
rect 363 220 364 222
rect 349 219 364 220
rect 372 222 376 223
rect 372 220 373 222
rect 375 220 376 222
rect 372 219 376 220
rect 499 222 563 223
rect 499 220 500 222
rect 502 220 560 222
rect 562 220 563 222
rect 499 219 563 220
rect -690 211 744 214
rect -690 209 739 211
rect 741 209 744 211
rect -690 207 -687 209
rect -685 207 -675 209
rect -673 207 -661 209
rect -659 207 -649 209
rect -647 207 -605 209
rect -603 207 -595 209
rect -593 207 -551 209
rect -549 207 -541 209
rect -539 207 -527 209
rect -525 207 -506 209
rect -504 207 -492 209
rect -490 207 -471 209
rect -469 207 -425 209
rect -423 207 -415 209
rect -413 207 -402 209
rect -400 207 -390 209
rect -388 207 -376 209
rect -374 207 -364 209
rect -362 207 -320 209
rect -318 207 -310 209
rect -308 207 -266 209
rect -264 207 -256 209
rect -254 207 -242 209
rect -240 207 -221 209
rect -219 207 -207 209
rect -205 207 -186 209
rect -184 207 -140 209
rect -138 207 -130 209
rect -128 207 -117 209
rect -115 207 -105 209
rect -103 207 -91 209
rect -89 207 -79 209
rect -77 207 -35 209
rect -33 207 -25 209
rect -23 207 19 209
rect 21 207 29 209
rect 31 207 43 209
rect 45 207 64 209
rect 66 207 78 209
rect 80 207 99 209
rect 101 207 145 209
rect 147 207 155 209
rect 157 207 168 209
rect 170 207 180 209
rect 182 207 194 209
rect 196 207 206 209
rect 208 207 250 209
rect 252 207 260 209
rect 262 207 304 209
rect 306 207 314 209
rect 316 207 328 209
rect 330 207 349 209
rect 351 207 363 209
rect 365 207 384 209
rect 386 207 430 209
rect 432 207 440 209
rect 442 207 457 209
rect 459 207 467 209
rect 469 207 517 209
rect 519 207 527 209
rect 529 207 583 209
rect 585 207 595 209
rect 597 207 744 209
rect -690 206 744 207
rect -682 185 -678 193
rect -674 192 -670 201
rect -672 190 -670 192
rect -690 183 -678 185
rect -690 181 -688 183
rect -686 181 -681 183
rect -679 181 -678 183
rect -690 179 -678 181
rect -674 186 -670 190
rect -674 184 -673 186
rect -671 184 -670 186
rect -656 185 -652 193
rect -648 192 -644 201
rect -646 190 -644 192
rect -674 174 -670 184
rect -664 183 -652 185
rect -664 181 -663 183
rect -661 181 -655 183
rect -653 181 -652 183
rect -664 179 -652 181
rect -648 186 -644 190
rect -648 184 -647 186
rect -645 184 -644 186
rect -672 172 -670 174
rect -674 169 -670 172
rect -648 174 -644 184
rect -635 192 -622 193
rect -635 190 -634 192
rect -632 190 -622 192
rect -635 187 -622 190
rect -618 190 -614 193
rect -618 188 -617 190
rect -615 188 -614 190
rect -594 193 -590 201
rect -592 191 -590 193
rect -635 183 -629 187
rect -635 181 -633 183
rect -631 181 -629 183
rect -635 180 -629 181
rect -618 184 -614 188
rect -618 183 -605 184
rect -618 181 -611 183
rect -609 181 -605 183
rect -618 180 -605 181
rect -646 172 -644 174
rect -635 175 -621 176
rect -635 173 -626 175
rect -624 174 -621 175
rect -619 174 -613 176
rect -624 173 -613 174
rect -635 172 -613 173
rect -594 185 -590 191
rect -594 183 -593 185
rect -591 183 -590 185
rect -648 169 -644 172
rect -682 167 -670 169
rect -682 165 -674 167
rect -672 165 -670 167
rect -682 163 -670 165
rect -656 167 -644 169
rect -656 165 -648 167
rect -646 165 -644 167
rect -656 163 -644 165
rect -627 164 -621 172
rect -594 172 -590 183
rect -581 192 -568 193
rect -581 190 -580 192
rect -578 190 -568 192
rect -581 187 -568 190
rect -564 190 -560 193
rect -564 188 -563 190
rect -561 188 -560 190
rect -540 193 -536 201
rect -519 200 -502 201
rect -519 198 -517 200
rect -515 198 -502 200
rect -519 197 -502 198
rect -514 195 -502 197
rect -538 191 -536 193
rect -581 183 -575 187
rect -581 181 -579 183
rect -577 181 -575 183
rect -581 180 -575 181
rect -564 184 -560 188
rect -564 183 -551 184
rect -564 181 -557 183
rect -555 181 -551 183
rect -564 180 -551 181
rect -581 175 -567 176
rect -581 173 -572 175
rect -570 174 -567 175
rect -565 174 -559 176
rect -570 173 -559 174
rect -581 172 -559 173
rect -540 185 -536 191
rect -522 187 -518 193
rect -540 183 -539 185
rect -537 183 -536 185
rect -592 170 -590 172
rect -594 168 -590 170
rect -603 165 -590 168
rect -603 164 -594 165
rect -595 163 -594 164
rect -592 163 -590 165
rect -595 155 -590 163
rect -573 164 -567 172
rect -540 172 -536 183
rect -530 186 -518 187
rect -530 184 -529 186
rect -527 184 -523 186
rect -521 184 -518 186
rect -506 191 -502 195
rect -484 200 -467 201
rect -484 198 -482 200
rect -480 198 -467 200
rect -484 197 -467 198
rect -479 195 -467 197
rect -471 193 -467 195
rect -506 189 -505 191
rect -503 189 -502 191
rect -530 183 -518 184
rect -514 183 -510 185
rect -530 179 -526 183
rect -514 181 -513 183
rect -511 181 -510 183
rect -514 179 -510 181
rect -538 170 -536 172
rect -522 178 -510 179
rect -522 176 -513 178
rect -511 176 -510 178
rect -522 175 -510 176
rect -522 171 -518 175
rect -540 168 -536 170
rect -549 165 -536 168
rect -506 167 -502 189
rect -487 187 -483 193
rect -495 186 -483 187
rect -495 184 -494 186
rect -492 184 -488 186
rect -486 184 -483 186
rect -471 191 -470 193
rect -468 191 -467 193
rect -495 183 -483 184
rect -479 183 -475 185
rect -495 179 -491 183
rect -479 181 -478 183
rect -476 181 -475 183
rect -479 179 -475 181
rect -487 178 -475 179
rect -487 176 -482 178
rect -480 176 -475 178
rect -487 175 -475 176
rect -487 171 -483 175
rect -471 167 -467 191
rect -455 192 -442 193
rect -455 190 -454 192
rect -452 190 -442 192
rect -455 187 -442 190
rect -438 191 -434 193
rect -438 189 -437 191
rect -435 189 -434 191
rect -414 193 -410 201
rect -412 191 -410 193
rect -414 189 -410 191
rect -455 183 -449 187
rect -455 181 -453 183
rect -451 181 -449 183
rect -455 180 -449 181
rect -438 184 -434 189
rect -438 183 -425 184
rect -438 181 -431 183
rect -429 181 -425 183
rect -438 180 -425 181
rect -455 175 -441 176
rect -455 173 -446 175
rect -444 174 -441 175
rect -439 174 -433 176
rect -444 173 -433 174
rect -455 172 -433 173
rect -414 187 -413 189
rect -411 187 -410 189
rect -549 164 -540 165
rect -541 163 -540 164
rect -538 163 -536 165
rect -541 155 -536 163
rect -511 166 -502 167
rect -511 164 -509 166
rect -507 164 -502 166
rect -511 163 -502 164
rect -476 166 -467 167
rect -476 164 -474 166
rect -472 164 -467 166
rect -476 163 -467 164
rect -511 159 -505 163
rect -511 157 -509 159
rect -507 157 -505 159
rect -511 156 -505 157
rect -476 159 -470 163
rect -476 157 -474 159
rect -472 157 -470 159
rect -476 156 -470 157
rect -447 164 -441 172
rect -414 172 -410 187
rect -397 185 -393 193
rect -389 192 -385 201
rect -387 190 -385 192
rect -405 183 -393 185
rect -405 181 -403 183
rect -401 181 -396 183
rect -394 181 -393 183
rect -405 179 -393 181
rect -389 186 -385 190
rect -389 184 -388 186
rect -386 184 -385 186
rect -371 185 -367 193
rect -363 192 -359 201
rect -361 190 -359 192
rect -412 170 -410 172
rect -414 168 -410 170
rect -389 174 -385 184
rect -379 183 -367 185
rect -379 181 -378 183
rect -376 181 -370 183
rect -368 181 -367 183
rect -379 179 -367 181
rect -363 186 -359 190
rect -363 184 -362 186
rect -360 184 -359 186
rect -387 172 -385 174
rect -389 169 -385 172
rect -363 174 -359 184
rect -350 192 -337 193
rect -350 190 -349 192
rect -347 190 -337 192
rect -350 187 -337 190
rect -333 190 -329 193
rect -333 188 -332 190
rect -330 188 -329 190
rect -309 193 -305 201
rect -307 191 -305 193
rect -350 183 -344 187
rect -350 181 -348 183
rect -346 181 -344 183
rect -350 180 -344 181
rect -333 184 -329 188
rect -333 183 -320 184
rect -333 181 -326 183
rect -324 181 -320 183
rect -333 180 -320 181
rect -361 172 -359 174
rect -350 175 -336 176
rect -350 173 -341 175
rect -339 174 -336 175
rect -334 174 -328 176
rect -339 173 -328 174
rect -350 172 -328 173
rect -309 185 -305 191
rect -309 183 -308 185
rect -306 183 -305 185
rect -363 169 -359 172
rect -423 165 -410 168
rect -423 164 -414 165
rect -415 163 -414 164
rect -412 163 -410 165
rect -397 167 -385 169
rect -397 165 -389 167
rect -387 165 -385 167
rect -397 163 -385 165
rect -371 167 -359 169
rect -371 165 -363 167
rect -361 165 -359 167
rect -371 163 -359 165
rect -471 150 -464 151
rect -415 155 -410 163
rect -342 164 -336 172
rect -309 172 -305 183
rect -296 192 -283 193
rect -296 190 -295 192
rect -293 190 -283 192
rect -296 187 -283 190
rect -279 190 -275 193
rect -279 188 -278 190
rect -276 188 -275 190
rect -255 193 -251 201
rect -234 200 -217 201
rect -234 198 -232 200
rect -230 198 -217 200
rect -234 197 -217 198
rect -229 195 -217 197
rect -253 191 -251 193
rect -296 183 -290 187
rect -296 181 -294 183
rect -292 181 -290 183
rect -296 180 -290 181
rect -279 184 -275 188
rect -279 183 -266 184
rect -279 181 -272 183
rect -270 181 -266 183
rect -279 180 -266 181
rect -296 175 -282 176
rect -296 173 -287 175
rect -285 174 -282 175
rect -280 174 -274 176
rect -285 173 -274 174
rect -296 172 -274 173
rect -255 185 -251 191
rect -237 187 -233 193
rect -255 183 -254 185
rect -252 183 -251 185
rect -307 170 -305 172
rect -309 168 -305 170
rect -318 165 -305 168
rect -318 164 -309 165
rect -310 163 -309 164
rect -307 163 -305 165
rect -310 155 -305 163
rect -288 164 -282 172
rect -255 172 -251 183
rect -245 186 -233 187
rect -245 184 -244 186
rect -242 184 -238 186
rect -236 184 -233 186
rect -221 191 -217 195
rect -199 200 -182 201
rect -199 198 -197 200
rect -195 198 -182 200
rect -199 197 -182 198
rect -194 195 -182 197
rect -186 193 -182 195
rect -221 189 -220 191
rect -218 189 -217 191
rect -245 183 -233 184
rect -229 183 -225 185
rect -245 179 -241 183
rect -229 181 -228 183
rect -226 181 -225 183
rect -229 179 -225 181
rect -253 170 -251 172
rect -237 178 -225 179
rect -237 176 -228 178
rect -226 176 -225 178
rect -237 175 -225 176
rect -237 171 -233 175
rect -255 168 -251 170
rect -264 165 -251 168
rect -221 167 -217 189
rect -202 187 -198 193
rect -210 186 -198 187
rect -210 184 -209 186
rect -207 184 -203 186
rect -201 184 -198 186
rect -186 191 -185 193
rect -183 191 -182 193
rect -210 183 -198 184
rect -194 183 -190 185
rect -210 179 -206 183
rect -194 181 -193 183
rect -191 181 -190 183
rect -194 179 -190 181
rect -202 178 -190 179
rect -202 176 -197 178
rect -195 176 -190 178
rect -202 175 -190 176
rect -202 171 -198 175
rect -186 167 -182 191
rect -170 192 -157 193
rect -170 190 -169 192
rect -167 190 -157 192
rect -170 187 -157 190
rect -153 191 -149 193
rect -153 189 -152 191
rect -150 189 -149 191
rect -129 193 -125 201
rect -127 191 -125 193
rect -129 189 -125 191
rect -170 183 -164 187
rect -170 181 -168 183
rect -166 181 -164 183
rect -170 180 -164 181
rect -153 184 -149 189
rect -153 183 -140 184
rect -153 181 -146 183
rect -144 181 -140 183
rect -153 180 -140 181
rect -170 175 -156 176
rect -170 173 -161 175
rect -159 174 -156 175
rect -154 174 -148 176
rect -159 173 -148 174
rect -170 172 -148 173
rect -129 187 -128 189
rect -126 187 -125 189
rect -264 164 -255 165
rect -256 163 -255 164
rect -253 163 -251 165
rect -256 155 -251 163
rect -226 166 -217 167
rect -226 164 -224 166
rect -222 164 -217 166
rect -226 163 -217 164
rect -191 166 -182 167
rect -191 164 -189 166
rect -187 164 -182 166
rect -191 163 -182 164
rect -226 159 -220 163
rect -226 157 -224 159
rect -222 157 -220 159
rect -226 156 -220 157
rect -191 159 -185 163
rect -191 157 -189 159
rect -187 157 -185 159
rect -191 156 -185 157
rect -162 164 -156 172
rect -129 172 -125 187
rect -112 185 -108 193
rect -104 192 -100 201
rect -102 190 -100 192
rect -120 183 -108 185
rect -120 181 -118 183
rect -116 181 -111 183
rect -109 181 -108 183
rect -120 179 -108 181
rect -104 186 -100 190
rect -104 184 -103 186
rect -101 184 -100 186
rect -86 185 -82 193
rect -78 192 -74 201
rect -76 190 -74 192
rect -127 170 -125 172
rect -129 168 -125 170
rect -104 174 -100 184
rect -94 183 -82 185
rect -94 181 -93 183
rect -91 181 -85 183
rect -83 181 -82 183
rect -94 179 -82 181
rect -78 186 -74 190
rect -78 184 -77 186
rect -75 184 -74 186
rect -102 172 -100 174
rect -104 169 -100 172
rect -78 174 -74 184
rect -65 192 -52 193
rect -65 190 -64 192
rect -62 190 -52 192
rect -65 187 -52 190
rect -48 190 -44 193
rect -48 188 -47 190
rect -45 188 -44 190
rect -24 193 -20 201
rect -22 191 -20 193
rect -65 183 -59 187
rect -65 181 -63 183
rect -61 181 -59 183
rect -65 180 -59 181
rect -48 184 -44 188
rect -48 183 -35 184
rect -48 181 -41 183
rect -39 181 -35 183
rect -48 180 -35 181
rect -76 172 -74 174
rect -65 175 -51 176
rect -65 173 -56 175
rect -54 174 -51 175
rect -49 174 -43 176
rect -54 173 -43 174
rect -65 172 -43 173
rect -24 185 -20 191
rect -24 183 -23 185
rect -21 183 -20 185
rect -78 169 -74 172
rect -138 165 -125 168
rect -138 164 -129 165
rect -130 163 -129 164
rect -127 163 -125 165
rect -112 167 -100 169
rect -112 165 -104 167
rect -102 165 -100 167
rect -112 163 -100 165
rect -86 167 -74 169
rect -86 165 -78 167
rect -76 165 -74 167
rect -86 163 -74 165
rect -186 150 -179 151
rect -130 155 -125 163
rect -57 164 -51 172
rect -24 172 -20 183
rect -11 192 2 193
rect -11 190 -10 192
rect -8 190 2 192
rect -11 187 2 190
rect 6 190 10 193
rect 6 188 7 190
rect 9 188 10 190
rect 30 193 34 201
rect 51 200 68 201
rect 51 198 53 200
rect 55 198 68 200
rect 51 197 68 198
rect 56 195 68 197
rect 32 191 34 193
rect -11 183 -5 187
rect -11 181 -9 183
rect -7 181 -5 183
rect -11 180 -5 181
rect 6 184 10 188
rect 6 183 19 184
rect 6 181 13 183
rect 15 181 19 183
rect 6 180 19 181
rect -11 175 3 176
rect -11 173 -2 175
rect 0 174 3 175
rect 5 174 11 176
rect 0 173 11 174
rect -11 172 11 173
rect 30 185 34 191
rect 48 187 52 193
rect 30 183 31 185
rect 33 183 34 185
rect -22 170 -20 172
rect -24 168 -20 170
rect -33 165 -20 168
rect -33 164 -24 165
rect -25 163 -24 164
rect -22 163 -20 165
rect -25 155 -20 163
rect -3 164 3 172
rect 30 172 34 183
rect 40 186 52 187
rect 40 184 41 186
rect 43 184 47 186
rect 49 184 52 186
rect 64 191 68 195
rect 86 200 103 201
rect 86 198 88 200
rect 90 198 103 200
rect 86 197 103 198
rect 91 195 103 197
rect 99 193 103 195
rect 64 189 65 191
rect 67 189 68 191
rect 40 183 52 184
rect 56 183 60 185
rect 40 179 44 183
rect 56 181 57 183
rect 59 181 60 183
rect 56 179 60 181
rect 32 170 34 172
rect 48 178 60 179
rect 48 176 57 178
rect 59 176 60 178
rect 48 175 60 176
rect 48 171 52 175
rect 30 168 34 170
rect 21 165 34 168
rect 64 167 68 189
rect 83 187 87 193
rect 75 186 87 187
rect 75 184 76 186
rect 78 184 82 186
rect 84 184 87 186
rect 99 191 100 193
rect 102 191 103 193
rect 75 183 87 184
rect 91 183 95 185
rect 75 179 79 183
rect 91 181 92 183
rect 94 181 95 183
rect 91 179 95 181
rect 83 178 95 179
rect 83 176 88 178
rect 90 176 95 178
rect 83 175 95 176
rect 83 171 87 175
rect 99 167 103 191
rect 115 192 128 193
rect 115 190 116 192
rect 118 190 128 192
rect 115 187 128 190
rect 132 191 136 193
rect 132 189 133 191
rect 135 189 136 191
rect 156 193 160 201
rect 158 191 160 193
rect 156 189 160 191
rect 115 183 121 187
rect 115 181 117 183
rect 119 181 121 183
rect 115 180 121 181
rect 132 184 136 189
rect 132 183 145 184
rect 132 181 139 183
rect 141 181 145 183
rect 132 180 145 181
rect 115 175 129 176
rect 115 173 124 175
rect 126 174 129 175
rect 131 174 137 176
rect 126 173 137 174
rect 115 172 137 173
rect 156 187 157 189
rect 159 187 160 189
rect 21 164 30 165
rect 29 163 30 164
rect 32 163 34 165
rect 29 155 34 163
rect 59 166 68 167
rect 59 164 61 166
rect 63 164 68 166
rect 59 163 68 164
rect 94 166 103 167
rect 94 164 96 166
rect 98 164 103 166
rect 94 163 103 164
rect 59 159 65 163
rect 59 157 61 159
rect 63 157 65 159
rect 59 156 65 157
rect 94 159 100 163
rect 94 157 96 159
rect 98 157 100 159
rect 94 156 100 157
rect 123 164 129 172
rect 156 172 160 187
rect 173 185 177 193
rect 181 192 185 201
rect 183 190 185 192
rect 165 183 177 185
rect 165 181 167 183
rect 169 181 174 183
rect 176 181 177 183
rect 165 179 177 181
rect 181 186 185 190
rect 181 184 182 186
rect 184 184 185 186
rect 199 185 203 193
rect 207 192 211 201
rect 209 190 211 192
rect 158 170 160 172
rect 156 168 160 170
rect 181 174 185 184
rect 191 183 203 185
rect 191 181 192 183
rect 194 181 200 183
rect 202 181 203 183
rect 191 179 203 181
rect 207 186 211 190
rect 207 184 208 186
rect 210 184 211 186
rect 183 172 185 174
rect 181 169 185 172
rect 207 174 211 184
rect 220 192 233 193
rect 220 190 221 192
rect 223 190 233 192
rect 220 187 233 190
rect 237 190 241 193
rect 237 188 238 190
rect 240 188 241 190
rect 261 193 265 201
rect 263 191 265 193
rect 220 183 226 187
rect 220 181 222 183
rect 224 181 226 183
rect 220 180 226 181
rect 237 184 241 188
rect 237 183 250 184
rect 237 181 244 183
rect 246 181 250 183
rect 237 180 250 181
rect 209 172 211 174
rect 220 175 234 176
rect 220 173 229 175
rect 231 174 234 175
rect 236 174 242 176
rect 231 173 242 174
rect 220 172 242 173
rect 261 185 265 191
rect 261 183 262 185
rect 264 183 265 185
rect 207 169 211 172
rect 147 165 160 168
rect 147 164 156 165
rect 155 163 156 164
rect 158 163 160 165
rect 173 167 185 169
rect 173 165 181 167
rect 183 165 185 167
rect 173 163 185 165
rect 199 167 211 169
rect 199 165 207 167
rect 209 165 211 167
rect 199 163 211 165
rect 99 150 106 151
rect 155 155 160 163
rect 228 164 234 172
rect 261 172 265 183
rect 274 192 287 193
rect 274 190 275 192
rect 277 190 287 192
rect 274 187 287 190
rect 291 190 295 193
rect 291 188 292 190
rect 294 188 295 190
rect 315 193 319 201
rect 336 200 353 201
rect 336 198 338 200
rect 340 198 353 200
rect 336 197 353 198
rect 341 195 353 197
rect 317 191 319 193
rect 274 183 280 187
rect 274 181 276 183
rect 278 181 280 183
rect 274 180 280 181
rect 291 184 295 188
rect 291 183 304 184
rect 291 181 298 183
rect 300 181 304 183
rect 291 180 304 181
rect 274 175 288 176
rect 274 173 283 175
rect 285 174 288 175
rect 290 174 296 176
rect 285 173 296 174
rect 274 172 296 173
rect 315 185 319 191
rect 333 187 337 193
rect 315 183 316 185
rect 318 183 319 185
rect 263 170 265 172
rect 261 168 265 170
rect 252 165 265 168
rect 252 164 261 165
rect 260 163 261 164
rect 263 163 265 165
rect 260 155 265 163
rect 282 164 288 172
rect 315 172 319 183
rect 325 186 337 187
rect 325 184 326 186
rect 328 184 332 186
rect 334 184 337 186
rect 349 191 353 195
rect 371 200 388 201
rect 371 198 373 200
rect 375 198 388 200
rect 371 197 388 198
rect 376 195 388 197
rect 384 193 388 195
rect 349 189 350 191
rect 352 189 353 191
rect 325 183 337 184
rect 341 183 345 185
rect 325 179 329 183
rect 341 181 342 183
rect 344 181 345 183
rect 341 179 345 181
rect 317 170 319 172
rect 333 178 345 179
rect 333 176 342 178
rect 344 176 345 178
rect 333 175 345 176
rect 333 171 337 175
rect 315 168 319 170
rect 306 165 319 168
rect 349 167 353 189
rect 368 187 372 193
rect 360 186 372 187
rect 360 184 361 186
rect 363 184 367 186
rect 369 184 372 186
rect 384 191 385 193
rect 387 191 388 193
rect 360 183 372 184
rect 376 183 380 185
rect 360 179 364 183
rect 376 181 377 183
rect 379 181 380 183
rect 376 179 380 181
rect 368 178 380 179
rect 368 176 373 178
rect 375 176 380 178
rect 368 175 380 176
rect 368 171 372 175
rect 384 167 388 191
rect 400 192 413 193
rect 400 190 401 192
rect 403 190 413 192
rect 400 187 413 190
rect 417 191 421 193
rect 417 189 418 191
rect 420 189 421 191
rect 441 193 445 201
rect 443 191 445 193
rect 441 189 445 191
rect 400 183 406 187
rect 400 181 402 183
rect 404 181 406 183
rect 400 180 406 181
rect 417 184 421 189
rect 417 183 430 184
rect 417 181 424 183
rect 426 181 430 183
rect 417 180 430 181
rect 400 175 414 176
rect 400 173 409 175
rect 411 174 414 175
rect 416 174 422 176
rect 411 173 422 174
rect 400 172 422 173
rect 441 187 442 189
rect 444 187 445 189
rect 306 164 315 165
rect 314 163 315 164
rect 317 163 319 165
rect 314 155 319 163
rect 344 166 353 167
rect 344 164 346 166
rect 348 164 353 166
rect 344 163 353 164
rect 379 166 388 167
rect 379 164 381 166
rect 383 164 388 166
rect 379 163 388 164
rect 344 159 350 163
rect 344 157 346 159
rect 348 157 350 159
rect 344 156 350 157
rect 379 159 385 163
rect 379 157 381 159
rect 383 157 385 159
rect 379 156 385 157
rect 408 164 414 172
rect 441 172 445 187
rect 443 170 445 172
rect 441 168 445 170
rect 432 165 445 168
rect 432 164 441 165
rect 440 163 441 164
rect 443 163 445 165
rect 384 150 391 151
rect 440 155 445 163
rect 454 193 458 201
rect 454 191 456 193
rect 454 187 458 191
rect 514 193 518 201
rect 580 199 584 201
rect 580 197 581 199
rect 583 197 584 199
rect 478 192 482 193
rect 478 190 479 192
rect 481 190 482 192
rect 454 185 455 187
rect 457 185 458 187
rect 454 172 458 185
rect 478 184 482 190
rect 486 190 500 193
rect 486 188 497 190
rect 499 188 500 190
rect 486 187 500 188
rect 514 191 516 193
rect 514 187 518 191
rect 538 192 542 193
rect 538 190 539 192
rect 541 190 542 192
rect 469 183 482 184
rect 469 181 473 183
rect 475 181 482 183
rect 469 180 482 181
rect 493 183 499 187
rect 493 181 495 183
rect 497 181 499 183
rect 493 180 499 181
rect 514 185 515 187
rect 517 185 518 187
rect 454 170 456 172
rect 454 168 458 170
rect 477 174 483 176
rect 485 175 499 176
rect 485 174 489 175
rect 477 173 489 174
rect 491 173 499 175
rect 477 172 499 173
rect 514 172 518 185
rect 538 184 542 190
rect 546 192 559 193
rect 546 190 551 192
rect 553 190 559 192
rect 546 187 559 190
rect 529 183 542 184
rect 529 181 533 183
rect 535 181 542 183
rect 529 180 542 181
rect 553 183 559 187
rect 553 181 555 183
rect 557 181 559 183
rect 553 180 559 181
rect 580 192 584 197
rect 580 190 582 192
rect 454 165 467 168
rect 454 163 456 165
rect 458 164 467 165
rect 458 163 459 164
rect 454 155 459 163
rect 485 164 491 172
rect 514 170 516 172
rect 514 168 518 170
rect 537 174 543 176
rect 545 175 563 176
rect 545 174 560 175
rect 537 173 560 174
rect 562 173 563 175
rect 537 172 563 173
rect 580 174 584 190
rect 588 185 592 193
rect 588 183 600 185
rect 588 181 589 183
rect 591 181 597 183
rect 599 181 600 183
rect 588 179 600 181
rect 580 172 582 174
rect 514 165 527 168
rect 514 163 516 165
rect 518 164 527 165
rect 518 163 519 164
rect 514 155 519 163
rect 545 164 551 172
rect 580 169 584 172
rect 580 167 592 169
rect 580 165 582 167
rect 584 165 592 167
rect 580 163 592 165
rect -738 149 604 150
rect -738 147 -687 149
rect -685 147 -675 149
rect -673 147 -661 149
rect -659 147 -649 149
rect -647 147 -639 149
rect -637 147 -625 149
rect -623 147 -585 149
rect -583 147 -571 149
rect -569 147 -459 149
rect -457 147 -445 149
rect -443 147 -402 149
rect -400 147 -390 149
rect -388 147 -376 149
rect -374 147 -364 149
rect -362 147 -354 149
rect -352 147 -340 149
rect -338 147 -300 149
rect -298 147 -286 149
rect -284 147 -174 149
rect -172 147 -160 149
rect -158 147 -117 149
rect -115 147 -105 149
rect -103 147 -91 149
rect -89 147 -79 149
rect -77 147 -69 149
rect -67 147 -55 149
rect -53 147 -15 149
rect -13 147 -1 149
rect 1 147 111 149
rect 113 147 125 149
rect 127 147 168 149
rect 170 147 180 149
rect 182 147 194 149
rect 196 147 206 149
rect 208 147 216 149
rect 218 147 230 149
rect 232 147 270 149
rect 272 147 284 149
rect 286 147 396 149
rect 398 147 410 149
rect 412 147 487 149
rect 489 147 501 149
rect 503 147 547 149
rect 549 147 561 149
rect 563 147 583 149
rect 585 147 595 149
rect 597 147 604 149
rect -738 143 604 147
rect -738 141 -733 143
rect -731 141 604 143
rect -738 137 604 141
rect -738 135 -687 137
rect -685 135 -675 137
rect -673 135 -661 137
rect -659 135 -649 137
rect -647 135 -639 137
rect -637 135 -625 137
rect -623 135 -585 137
rect -583 135 -571 137
rect -569 135 -459 137
rect -457 135 -445 137
rect -443 135 -402 137
rect -400 135 -390 137
rect -388 135 -376 137
rect -374 135 -364 137
rect -362 135 -354 137
rect -352 135 -340 137
rect -338 135 -300 137
rect -298 135 -286 137
rect -284 135 -174 137
rect -172 135 -160 137
rect -158 135 -117 137
rect -115 135 -105 137
rect -103 135 -91 137
rect -89 135 -79 137
rect -77 135 -69 137
rect -67 135 -55 137
rect -53 135 -15 137
rect -13 135 -1 137
rect 1 135 111 137
rect 113 135 125 137
rect 127 135 168 137
rect 170 135 180 137
rect 182 135 194 137
rect 196 135 206 137
rect 208 135 216 137
rect 218 135 230 137
rect 232 135 270 137
rect 272 135 284 137
rect 286 135 396 137
rect 398 135 410 137
rect 412 135 487 137
rect 489 135 501 137
rect 503 135 547 137
rect 549 135 561 137
rect 563 135 583 137
rect 585 135 595 137
rect 597 135 604 137
rect -738 134 604 135
rect -682 119 -670 121
rect -682 117 -674 119
rect -672 117 -670 119
rect -682 115 -670 117
rect -656 119 -644 121
rect -656 117 -648 119
rect -646 117 -644 119
rect -656 115 -644 117
rect -674 112 -670 115
rect -672 110 -670 112
rect -690 103 -678 105
rect -690 101 -688 103
rect -686 101 -681 103
rect -679 101 -678 103
rect -690 99 -678 101
rect -682 91 -678 99
rect -674 100 -670 110
rect -648 112 -644 115
rect -627 112 -621 120
rect -595 121 -590 129
rect -595 120 -594 121
rect -603 119 -594 120
rect -592 119 -590 121
rect -603 116 -590 119
rect -646 110 -644 112
rect -674 98 -673 100
rect -671 98 -670 100
rect -664 103 -652 105
rect -664 101 -663 103
rect -661 101 -655 103
rect -653 101 -652 103
rect -664 99 -652 101
rect -674 94 -670 98
rect -672 92 -670 94
rect -674 83 -670 92
rect -656 91 -652 99
rect -648 100 -644 110
rect -635 111 -613 112
rect -635 109 -626 111
rect -624 110 -613 111
rect -624 109 -621 110
rect -635 108 -621 109
rect -619 108 -613 110
rect -594 114 -590 116
rect -592 112 -590 114
rect -573 112 -567 120
rect -541 121 -536 129
rect -471 133 -453 134
rect -511 127 -505 128
rect -511 125 -509 127
rect -507 125 -505 127
rect -541 120 -540 121
rect -549 119 -540 120
rect -538 119 -536 121
rect -549 116 -536 119
rect -511 121 -505 125
rect -476 127 -470 128
rect -476 125 -474 127
rect -472 125 -470 127
rect -476 121 -470 125
rect -511 120 -502 121
rect -511 118 -509 120
rect -507 118 -502 120
rect -511 117 -502 118
rect -476 120 -467 121
rect -476 118 -474 120
rect -472 118 -467 120
rect -476 117 -467 118
rect -648 98 -647 100
rect -645 98 -644 100
rect -648 94 -644 98
rect -646 92 -644 94
rect -648 83 -644 92
rect -635 103 -629 104
rect -635 101 -633 103
rect -631 101 -629 103
rect -635 97 -629 101
rect -618 103 -605 104
rect -618 101 -611 103
rect -609 101 -605 103
rect -618 100 -605 101
rect -635 94 -622 97
rect -635 92 -634 94
rect -632 92 -622 94
rect -635 91 -622 92
rect -618 96 -614 100
rect -618 94 -617 96
rect -615 94 -614 96
rect -594 101 -590 112
rect -581 111 -559 112
rect -581 109 -572 111
rect -570 110 -559 111
rect -570 109 -567 110
rect -581 108 -567 109
rect -565 108 -559 110
rect -540 114 -536 116
rect -538 112 -536 114
rect -594 99 -593 101
rect -591 99 -590 101
rect -618 91 -614 94
rect -594 93 -590 99
rect -592 91 -590 93
rect -581 103 -575 104
rect -581 101 -579 103
rect -577 101 -575 103
rect -581 97 -575 101
rect -564 103 -551 104
rect -564 101 -557 103
rect -555 101 -551 103
rect -564 100 -551 101
rect -581 94 -568 97
rect -581 92 -580 94
rect -578 92 -568 94
rect -581 91 -568 92
rect -564 96 -560 100
rect -564 94 -563 96
rect -561 94 -560 96
rect -540 101 -536 112
rect -522 109 -518 113
rect -522 108 -510 109
rect -522 106 -513 108
rect -511 106 -510 108
rect -522 105 -510 106
rect -540 99 -539 101
rect -537 99 -536 101
rect -564 91 -560 94
rect -594 83 -590 91
rect -540 93 -536 99
rect -530 101 -526 105
rect -514 103 -510 105
rect -514 101 -513 103
rect -511 101 -510 103
rect -530 100 -518 101
rect -530 98 -529 100
rect -527 98 -523 100
rect -521 98 -518 100
rect -514 99 -510 101
rect -530 97 -518 98
rect -538 91 -536 93
rect -522 91 -518 97
rect -506 95 -502 117
rect -487 109 -483 113
rect -487 108 -475 109
rect -487 106 -482 108
rect -480 106 -475 108
rect -487 105 -475 106
rect -495 101 -491 105
rect -479 103 -475 105
rect -479 101 -478 103
rect -476 101 -475 103
rect -495 100 -483 101
rect -495 98 -494 100
rect -492 98 -488 100
rect -486 98 -483 100
rect -479 99 -475 101
rect -495 97 -483 98
rect -506 93 -505 95
rect -503 93 -502 95
rect -540 83 -536 91
rect -506 89 -502 93
rect -487 91 -483 97
rect -471 93 -467 117
rect -447 112 -441 120
rect -415 121 -410 129
rect -415 120 -414 121
rect -423 119 -414 120
rect -412 119 -410 121
rect -423 116 -410 119
rect -455 111 -433 112
rect -455 109 -446 111
rect -444 110 -433 111
rect -444 109 -441 110
rect -455 108 -441 109
rect -439 108 -433 110
rect -414 114 -410 116
rect -397 119 -385 121
rect -397 117 -389 119
rect -387 117 -385 119
rect -397 115 -385 117
rect -371 119 -359 121
rect -371 117 -363 119
rect -361 117 -359 119
rect -371 115 -359 117
rect -412 112 -410 114
rect -471 91 -470 93
rect -468 91 -467 93
rect -455 103 -449 104
rect -455 101 -453 103
rect -451 101 -449 103
rect -455 97 -449 101
rect -438 103 -425 104
rect -438 101 -431 103
rect -429 101 -425 103
rect -438 100 -425 101
rect -455 94 -442 97
rect -455 92 -454 94
rect -452 92 -442 94
rect -455 91 -442 92
rect -438 95 -434 100
rect -414 97 -410 112
rect -389 112 -385 115
rect -387 110 -385 112
rect -405 103 -393 105
rect -405 101 -403 103
rect -401 101 -396 103
rect -394 101 -393 103
rect -405 99 -393 101
rect -414 95 -413 97
rect -411 95 -410 97
rect -438 93 -437 95
rect -435 93 -434 95
rect -438 91 -434 93
rect -514 87 -502 89
rect -519 86 -502 87
rect -519 84 -517 86
rect -515 84 -502 86
rect -519 83 -502 84
rect -471 89 -467 91
rect -479 87 -467 89
rect -414 93 -410 95
rect -412 91 -410 93
rect -484 86 -467 87
rect -484 84 -482 86
rect -480 84 -467 86
rect -484 83 -467 84
rect -414 83 -410 91
rect -397 91 -393 99
rect -389 100 -385 110
rect -363 112 -359 115
rect -342 112 -336 120
rect -310 121 -305 129
rect -310 120 -309 121
rect -318 119 -309 120
rect -307 119 -305 121
rect -318 116 -305 119
rect -361 110 -359 112
rect -389 98 -388 100
rect -386 98 -385 100
rect -379 103 -367 105
rect -379 101 -378 103
rect -376 101 -370 103
rect -368 101 -367 103
rect -379 99 -367 101
rect -389 94 -385 98
rect -387 92 -385 94
rect -389 83 -385 92
rect -371 91 -367 99
rect -363 100 -359 110
rect -350 111 -328 112
rect -350 109 -341 111
rect -339 110 -328 111
rect -339 109 -336 110
rect -350 108 -336 109
rect -334 108 -328 110
rect -309 114 -305 116
rect -307 112 -305 114
rect -288 112 -282 120
rect -256 121 -251 129
rect -226 127 -220 128
rect -226 125 -224 127
rect -222 125 -220 127
rect -256 120 -255 121
rect -264 119 -255 120
rect -253 119 -251 121
rect -264 116 -251 119
rect -226 121 -220 125
rect -191 127 -185 128
rect -191 125 -189 127
rect -187 125 -185 127
rect -191 121 -185 125
rect -226 120 -217 121
rect -226 118 -224 120
rect -222 118 -217 120
rect -226 117 -217 118
rect -191 120 -182 121
rect -191 118 -189 120
rect -187 118 -182 120
rect -191 117 -182 118
rect -363 98 -362 100
rect -360 98 -359 100
rect -363 94 -359 98
rect -361 92 -359 94
rect -363 83 -359 92
rect -350 103 -344 104
rect -350 101 -348 103
rect -346 101 -344 103
rect -350 97 -344 101
rect -333 103 -320 104
rect -333 101 -326 103
rect -324 101 -320 103
rect -333 100 -320 101
rect -350 94 -337 97
rect -350 92 -349 94
rect -347 92 -337 94
rect -350 91 -337 92
rect -333 96 -329 100
rect -333 94 -332 96
rect -330 94 -329 96
rect -309 101 -305 112
rect -296 111 -274 112
rect -296 109 -287 111
rect -285 110 -274 111
rect -285 109 -282 110
rect -296 108 -282 109
rect -280 108 -274 110
rect -255 114 -251 116
rect -253 112 -251 114
rect -309 99 -308 101
rect -306 99 -305 101
rect -333 91 -329 94
rect -309 93 -305 99
rect -307 91 -305 93
rect -296 103 -290 104
rect -296 101 -294 103
rect -292 101 -290 103
rect -296 97 -290 101
rect -279 103 -266 104
rect -279 101 -272 103
rect -270 101 -266 103
rect -279 100 -266 101
rect -296 94 -283 97
rect -296 92 -295 94
rect -293 92 -283 94
rect -296 91 -283 92
rect -279 96 -275 100
rect -279 94 -278 96
rect -276 94 -275 96
rect -255 101 -251 112
rect -237 109 -233 113
rect -237 108 -225 109
rect -237 106 -228 108
rect -226 106 -225 108
rect -237 105 -225 106
rect -255 99 -254 101
rect -252 99 -251 101
rect -279 91 -275 94
rect -309 83 -305 91
rect -255 93 -251 99
rect -245 101 -241 105
rect -229 103 -225 105
rect -229 101 -228 103
rect -226 101 -225 103
rect -245 100 -233 101
rect -245 98 -244 100
rect -242 98 -238 100
rect -236 98 -233 100
rect -229 99 -225 101
rect -245 97 -233 98
rect -253 91 -251 93
rect -237 91 -233 97
rect -221 95 -217 117
rect -202 109 -198 113
rect -202 108 -190 109
rect -202 106 -197 108
rect -195 106 -190 108
rect -202 105 -190 106
rect -210 101 -206 105
rect -194 103 -190 105
rect -194 101 -193 103
rect -191 101 -190 103
rect -210 100 -198 101
rect -210 98 -209 100
rect -207 98 -203 100
rect -201 98 -198 100
rect -194 99 -190 101
rect -210 97 -198 98
rect -221 93 -220 95
rect -218 93 -217 95
rect -255 83 -251 91
rect -221 89 -217 93
rect -202 91 -198 97
rect -186 93 -182 117
rect -162 112 -156 120
rect -130 121 -125 129
rect -130 120 -129 121
rect -138 119 -129 120
rect -127 119 -125 121
rect -138 116 -125 119
rect -170 111 -148 112
rect -170 109 -161 111
rect -159 110 -148 111
rect -159 109 -156 110
rect -170 108 -156 109
rect -154 108 -148 110
rect -129 114 -125 116
rect -112 119 -100 121
rect -112 117 -104 119
rect -102 117 -100 119
rect -112 115 -100 117
rect -86 119 -74 121
rect -86 117 -78 119
rect -76 117 -74 119
rect -86 115 -74 117
rect -127 112 -125 114
rect -186 91 -185 93
rect -183 91 -182 93
rect -170 103 -164 104
rect -170 101 -168 103
rect -166 101 -164 103
rect -170 97 -164 101
rect -153 103 -140 104
rect -153 101 -146 103
rect -144 101 -140 103
rect -153 100 -140 101
rect -170 94 -157 97
rect -170 92 -169 94
rect -167 92 -157 94
rect -170 91 -157 92
rect -153 95 -149 100
rect -129 97 -125 112
rect -104 112 -100 115
rect -102 110 -100 112
rect -120 103 -108 105
rect -120 101 -118 103
rect -116 101 -111 103
rect -109 101 -108 103
rect -120 99 -108 101
rect -129 95 -128 97
rect -126 95 -125 97
rect -153 93 -152 95
rect -150 93 -149 95
rect -153 91 -149 93
rect -229 87 -217 89
rect -234 86 -217 87
rect -234 84 -232 86
rect -230 84 -217 86
rect -234 83 -217 84
rect -186 89 -182 91
rect -194 87 -182 89
rect -129 93 -125 95
rect -127 91 -125 93
rect -199 86 -182 87
rect -199 84 -197 86
rect -195 84 -182 86
rect -199 83 -182 84
rect -129 83 -125 91
rect -112 91 -108 99
rect -104 100 -100 110
rect -78 112 -74 115
rect -57 112 -51 120
rect -25 121 -20 129
rect -25 120 -24 121
rect -33 119 -24 120
rect -22 119 -20 121
rect -33 116 -20 119
rect -76 110 -74 112
rect -104 98 -103 100
rect -101 98 -100 100
rect -94 103 -82 105
rect -94 101 -93 103
rect -91 101 -85 103
rect -83 101 -82 103
rect -94 99 -82 101
rect -104 94 -100 98
rect -102 92 -100 94
rect -104 83 -100 92
rect -86 91 -82 99
rect -78 100 -74 110
rect -65 111 -43 112
rect -65 109 -56 111
rect -54 110 -43 111
rect -54 109 -51 110
rect -65 108 -51 109
rect -49 108 -43 110
rect -24 114 -20 116
rect -22 112 -20 114
rect -3 112 3 120
rect 29 121 34 129
rect 59 127 65 128
rect 59 125 61 127
rect 63 125 65 127
rect 29 120 30 121
rect 21 119 30 120
rect 32 119 34 121
rect 21 116 34 119
rect 59 121 65 125
rect 94 127 100 128
rect 94 125 96 127
rect 98 125 100 127
rect 94 121 100 125
rect 59 120 68 121
rect 59 118 61 120
rect 63 118 68 120
rect 59 117 68 118
rect 94 120 103 121
rect 94 118 96 120
rect 98 118 103 120
rect 94 117 103 118
rect -78 98 -77 100
rect -75 98 -74 100
rect -78 94 -74 98
rect -76 92 -74 94
rect -78 83 -74 92
rect -65 103 -59 104
rect -65 101 -63 103
rect -61 101 -59 103
rect -65 97 -59 101
rect -48 103 -35 104
rect -48 101 -41 103
rect -39 101 -35 103
rect -48 100 -35 101
rect -65 94 -52 97
rect -65 92 -64 94
rect -62 92 -52 94
rect -65 91 -52 92
rect -48 96 -44 100
rect -48 94 -47 96
rect -45 94 -44 96
rect -24 101 -20 112
rect -11 111 11 112
rect -11 109 -2 111
rect 0 110 11 111
rect 0 109 3 110
rect -11 108 3 109
rect 5 108 11 110
rect 30 114 34 116
rect 32 112 34 114
rect -24 99 -23 101
rect -21 99 -20 101
rect -48 91 -44 94
rect -24 93 -20 99
rect -22 91 -20 93
rect -11 103 -5 104
rect -11 101 -9 103
rect -7 101 -5 103
rect -11 97 -5 101
rect 6 103 19 104
rect 6 101 13 103
rect 15 101 19 103
rect 6 100 19 101
rect -11 94 2 97
rect -11 92 -10 94
rect -8 92 2 94
rect -11 91 2 92
rect 6 96 10 100
rect 6 94 7 96
rect 9 94 10 96
rect 30 101 34 112
rect 48 109 52 113
rect 48 108 60 109
rect 48 106 57 108
rect 59 106 60 108
rect 48 105 60 106
rect 30 99 31 101
rect 33 99 34 101
rect 6 91 10 94
rect -24 83 -20 91
rect 30 93 34 99
rect 40 101 44 105
rect 56 103 60 105
rect 56 101 57 103
rect 59 101 60 103
rect 40 100 52 101
rect 40 98 41 100
rect 43 98 47 100
rect 49 98 52 100
rect 56 99 60 101
rect 40 97 52 98
rect 32 91 34 93
rect 48 91 52 97
rect 64 95 68 117
rect 83 109 87 113
rect 83 108 95 109
rect 83 106 88 108
rect 90 106 95 108
rect 83 105 95 106
rect 75 101 79 105
rect 91 103 95 105
rect 91 101 92 103
rect 94 101 95 103
rect 75 100 87 101
rect 75 98 76 100
rect 78 98 82 100
rect 84 98 87 100
rect 91 99 95 101
rect 75 97 87 98
rect 64 93 65 95
rect 67 93 68 95
rect 30 83 34 91
rect 64 89 68 93
rect 83 91 87 97
rect 99 93 103 117
rect 123 112 129 120
rect 155 121 160 129
rect 155 120 156 121
rect 147 119 156 120
rect 158 119 160 121
rect 147 116 160 119
rect 115 111 137 112
rect 115 109 124 111
rect 126 110 137 111
rect 126 109 129 110
rect 115 108 129 109
rect 131 108 137 110
rect 156 114 160 116
rect 173 119 185 121
rect 173 117 181 119
rect 183 117 185 119
rect 173 115 185 117
rect 199 119 211 121
rect 199 117 207 119
rect 209 117 211 119
rect 199 115 211 117
rect 158 112 160 114
rect 99 91 100 93
rect 102 91 103 93
rect 115 103 121 104
rect 115 101 117 103
rect 119 101 121 103
rect 115 97 121 101
rect 132 103 145 104
rect 132 101 139 103
rect 141 101 145 103
rect 132 100 145 101
rect 115 94 128 97
rect 115 92 116 94
rect 118 92 128 94
rect 115 91 128 92
rect 132 95 136 100
rect 156 97 160 112
rect 181 112 185 115
rect 183 110 185 112
rect 165 103 177 105
rect 165 101 167 103
rect 169 101 174 103
rect 176 101 177 103
rect 165 99 177 101
rect 156 95 157 97
rect 159 95 160 97
rect 132 93 133 95
rect 135 93 136 95
rect 132 91 136 93
rect 56 87 68 89
rect 51 86 68 87
rect 51 84 53 86
rect 55 84 68 86
rect 51 83 68 84
rect 99 89 103 91
rect 91 87 103 89
rect 156 93 160 95
rect 158 91 160 93
rect 86 86 103 87
rect 86 84 88 86
rect 90 84 103 86
rect 86 83 103 84
rect 156 83 160 91
rect 173 91 177 99
rect 181 100 185 110
rect 207 112 211 115
rect 228 112 234 120
rect 260 121 265 129
rect 260 120 261 121
rect 252 119 261 120
rect 263 119 265 121
rect 252 116 265 119
rect 209 110 211 112
rect 181 98 182 100
rect 184 98 185 100
rect 191 103 203 105
rect 191 101 192 103
rect 194 101 200 103
rect 202 101 203 103
rect 191 99 203 101
rect 181 94 185 98
rect 183 92 185 94
rect 181 83 185 92
rect 199 91 203 99
rect 207 100 211 110
rect 220 111 242 112
rect 220 109 229 111
rect 231 110 242 111
rect 231 109 234 110
rect 220 108 234 109
rect 236 108 242 110
rect 261 114 265 116
rect 263 112 265 114
rect 282 112 288 120
rect 314 121 319 129
rect 344 127 350 128
rect 344 125 346 127
rect 348 125 350 127
rect 314 120 315 121
rect 306 119 315 120
rect 317 119 319 121
rect 306 116 319 119
rect 344 121 350 125
rect 379 127 385 128
rect 379 125 381 127
rect 383 125 385 127
rect 379 121 385 125
rect 344 120 353 121
rect 344 118 346 120
rect 348 118 353 120
rect 344 117 353 118
rect 379 120 388 121
rect 379 118 381 120
rect 383 118 388 120
rect 379 117 388 118
rect 207 98 208 100
rect 210 98 211 100
rect 207 94 211 98
rect 209 92 211 94
rect 207 83 211 92
rect 220 103 226 104
rect 220 101 222 103
rect 224 101 226 103
rect 220 97 226 101
rect 237 103 250 104
rect 237 101 244 103
rect 246 101 250 103
rect 237 100 250 101
rect 220 94 233 97
rect 220 92 221 94
rect 223 92 233 94
rect 220 91 233 92
rect 237 96 241 100
rect 237 94 238 96
rect 240 94 241 96
rect 261 101 265 112
rect 274 111 296 112
rect 274 109 283 111
rect 285 110 296 111
rect 285 109 288 110
rect 274 108 288 109
rect 290 108 296 110
rect 315 114 319 116
rect 317 112 319 114
rect 261 99 262 101
rect 264 99 265 101
rect 237 91 241 94
rect 261 93 265 99
rect 263 91 265 93
rect 274 103 280 104
rect 274 101 276 103
rect 278 101 280 103
rect 274 97 280 101
rect 291 103 304 104
rect 291 101 298 103
rect 300 101 304 103
rect 291 100 304 101
rect 274 94 287 97
rect 274 92 275 94
rect 277 92 287 94
rect 274 91 287 92
rect 291 96 295 100
rect 291 94 292 96
rect 294 94 295 96
rect 315 101 319 112
rect 333 109 337 113
rect 333 108 345 109
rect 333 106 342 108
rect 344 106 345 108
rect 333 105 345 106
rect 315 99 316 101
rect 318 99 319 101
rect 291 91 295 94
rect 261 83 265 91
rect 315 93 319 99
rect 325 101 329 105
rect 341 103 345 105
rect 341 101 342 103
rect 344 101 345 103
rect 325 100 337 101
rect 325 98 326 100
rect 328 98 332 100
rect 334 98 337 100
rect 341 99 345 101
rect 325 97 337 98
rect 317 91 319 93
rect 333 91 337 97
rect 349 95 353 117
rect 368 109 372 113
rect 368 108 380 109
rect 368 106 373 108
rect 375 106 380 108
rect 368 105 380 106
rect 360 101 364 105
rect 376 103 380 105
rect 376 101 377 103
rect 379 101 380 103
rect 360 100 372 101
rect 360 98 361 100
rect 363 98 367 100
rect 369 98 372 100
rect 376 99 380 101
rect 360 97 372 98
rect 349 93 350 95
rect 352 93 353 95
rect 315 83 319 91
rect 349 89 353 93
rect 368 91 372 97
rect 384 93 388 117
rect 408 112 414 120
rect 440 121 445 129
rect 440 120 441 121
rect 432 119 441 120
rect 443 119 445 121
rect 432 116 445 119
rect 400 111 422 112
rect 400 109 409 111
rect 411 110 422 111
rect 411 109 414 110
rect 400 108 414 109
rect 416 108 422 110
rect 441 114 445 116
rect 443 112 445 114
rect 384 91 385 93
rect 387 91 388 93
rect 400 103 406 104
rect 400 101 402 103
rect 404 101 406 103
rect 400 97 406 101
rect 417 103 430 104
rect 417 101 424 103
rect 426 101 430 103
rect 417 100 430 101
rect 400 94 413 97
rect 400 92 401 94
rect 403 92 413 94
rect 400 91 413 92
rect 417 95 421 100
rect 441 97 445 112
rect 441 95 442 97
rect 444 95 445 97
rect 417 93 418 95
rect 420 93 421 95
rect 417 91 421 93
rect 341 87 353 89
rect 336 86 353 87
rect 336 84 338 86
rect 340 84 353 86
rect 336 83 353 84
rect 384 89 388 91
rect 376 87 388 89
rect 441 93 445 95
rect 443 91 445 93
rect 371 86 388 87
rect 371 84 373 86
rect 375 84 388 86
rect 371 83 388 84
rect 441 83 445 91
rect 454 121 459 129
rect 454 119 456 121
rect 458 120 459 121
rect 458 119 467 120
rect 454 116 467 119
rect 454 114 458 116
rect 454 112 456 114
rect 454 101 458 112
rect 485 112 491 120
rect 514 121 519 129
rect 514 119 516 121
rect 518 120 519 121
rect 518 119 527 120
rect 514 116 527 119
rect 514 114 518 116
rect 514 112 516 114
rect 454 99 455 101
rect 457 99 458 101
rect 454 93 458 99
rect 477 111 499 112
rect 477 110 489 111
rect 477 108 483 110
rect 485 109 489 110
rect 491 109 499 111
rect 485 108 499 109
rect 469 103 482 104
rect 469 101 473 103
rect 475 101 482 103
rect 469 100 482 101
rect 454 91 456 93
rect 454 83 458 91
rect 478 94 482 100
rect 493 103 499 104
rect 493 101 495 103
rect 497 101 499 103
rect 493 97 499 101
rect 514 101 518 112
rect 545 112 551 120
rect 580 119 592 121
rect 580 117 582 119
rect 584 117 592 119
rect 580 115 592 117
rect 580 112 584 115
rect 514 99 515 101
rect 517 99 518 101
rect 478 92 479 94
rect 481 92 482 94
rect 478 91 482 92
rect 486 96 500 97
rect 486 94 497 96
rect 499 94 500 96
rect 486 91 500 94
rect 514 93 518 99
rect 537 111 559 112
rect 537 110 549 111
rect 537 108 543 110
rect 545 109 549 110
rect 551 109 559 111
rect 545 108 559 109
rect 580 110 582 112
rect 529 103 542 104
rect 529 101 533 103
rect 535 101 542 103
rect 529 100 542 101
rect 514 91 516 93
rect 514 83 518 91
rect 538 94 542 100
rect 553 103 559 104
rect 553 101 555 103
rect 557 101 559 103
rect 553 97 559 101
rect 538 92 539 94
rect 541 92 542 94
rect 538 91 542 92
rect 546 96 560 97
rect 546 94 557 96
rect 559 94 560 96
rect 546 91 560 94
rect 580 94 584 110
rect 588 103 600 105
rect 588 101 589 103
rect 591 101 597 103
rect 599 101 600 103
rect 588 99 600 101
rect 580 92 582 94
rect 580 87 584 92
rect 588 91 592 99
rect 580 85 581 87
rect 583 85 584 87
rect 580 83 584 85
rect -690 77 744 78
rect -690 75 -687 77
rect -685 75 -675 77
rect -673 75 -661 77
rect -659 75 -649 77
rect -647 75 -605 77
rect -603 75 -595 77
rect -593 75 -551 77
rect -549 75 -541 77
rect -539 75 -527 77
rect -525 75 -506 77
rect -504 75 -492 77
rect -490 75 -471 77
rect -469 75 -425 77
rect -423 75 -415 77
rect -413 75 -402 77
rect -400 75 -390 77
rect -388 75 -376 77
rect -374 75 -364 77
rect -362 75 -320 77
rect -318 75 -310 77
rect -308 75 -266 77
rect -264 75 -256 77
rect -254 75 -242 77
rect -240 75 -221 77
rect -219 75 -207 77
rect -205 75 -186 77
rect -184 75 -140 77
rect -138 75 -130 77
rect -128 75 -117 77
rect -115 75 -105 77
rect -103 75 -91 77
rect -89 75 -79 77
rect -77 75 -35 77
rect -33 75 -25 77
rect -23 75 19 77
rect 21 75 29 77
rect 31 75 43 77
rect 45 75 64 77
rect 66 75 78 77
rect 80 75 99 77
rect 101 75 145 77
rect 147 75 155 77
rect 157 75 168 77
rect 170 75 180 77
rect 182 75 194 77
rect 196 75 206 77
rect 208 75 250 77
rect 252 75 260 77
rect 262 75 304 77
rect 306 75 314 77
rect 316 75 328 77
rect 330 75 349 77
rect 351 75 363 77
rect 365 75 384 77
rect 386 75 430 77
rect 432 75 440 77
rect 442 75 457 77
rect 459 75 467 77
rect 469 75 517 77
rect 519 75 527 77
rect 529 75 583 77
rect 585 75 595 77
rect 597 75 744 77
rect -690 73 740 75
rect 742 73 744 75
rect -690 70 744 73
rect -674 64 -631 65
rect -674 62 -673 64
rect -671 62 -634 64
rect -632 62 -631 64
rect -674 61 -631 62
rect -540 64 -526 65
rect -540 62 -539 64
rect -537 62 -529 64
rect -527 62 -526 64
rect -540 61 -526 62
rect -506 64 -491 65
rect -506 62 -505 64
rect -503 62 -494 64
rect -492 62 -491 64
rect -506 61 -491 62
rect -483 64 -479 65
rect -483 62 -482 64
rect -480 62 -479 64
rect -483 61 -479 62
rect -389 64 -346 65
rect -389 62 -388 64
rect -386 62 -349 64
rect -347 62 -346 64
rect -389 61 -346 62
rect -255 64 -241 65
rect -255 62 -254 64
rect -252 62 -244 64
rect -242 62 -241 64
rect -255 61 -241 62
rect -221 64 -206 65
rect -221 62 -220 64
rect -218 62 -209 64
rect -207 62 -206 64
rect -221 61 -206 62
rect -198 64 -194 65
rect -198 62 -197 64
rect -195 62 -194 64
rect -198 61 -194 62
rect -104 64 -61 65
rect -104 62 -103 64
rect -101 62 -64 64
rect -62 62 -61 64
rect -104 61 -61 62
rect 30 64 44 65
rect 30 62 31 64
rect 33 62 41 64
rect 43 62 44 64
rect 30 61 44 62
rect 64 64 79 65
rect 64 62 65 64
rect 67 62 76 64
rect 78 62 79 64
rect 64 61 79 62
rect 87 64 91 65
rect 87 62 88 64
rect 90 62 91 64
rect 87 61 91 62
rect 181 64 224 65
rect 181 62 182 64
rect 184 62 221 64
rect 223 62 224 64
rect 181 61 224 62
rect 315 64 329 65
rect 315 62 316 64
rect 318 62 326 64
rect 328 62 329 64
rect 315 61 329 62
rect 349 64 364 65
rect 349 62 350 64
rect 352 62 361 64
rect 363 62 364 64
rect 349 61 364 62
rect 372 64 376 65
rect 372 62 373 64
rect 375 62 376 64
rect 372 61 376 62
rect 499 64 563 65
rect 499 62 500 64
rect 502 62 560 64
rect 562 62 563 64
rect 499 61 563 62
rect -689 56 -577 57
rect -689 54 -688 56
rect -686 54 -580 56
rect -578 54 -577 56
rect -689 53 -577 54
rect -514 56 -451 57
rect -514 54 -513 56
rect -511 54 -470 56
rect -468 54 -454 56
rect -452 54 -451 56
rect -514 53 -451 54
rect -404 56 -292 57
rect -404 54 -403 56
rect -401 54 -295 56
rect -293 54 -292 56
rect -404 53 -292 54
rect -229 56 -166 57
rect -229 54 -228 56
rect -226 54 -185 56
rect -183 54 -169 56
rect -167 54 -166 56
rect -229 53 -166 54
rect -119 56 -7 57
rect -119 54 -118 56
rect -116 54 -10 56
rect -8 54 -7 56
rect -119 53 -7 54
rect 56 56 119 57
rect 56 54 57 56
rect 59 54 100 56
rect 102 54 116 56
rect 118 54 119 56
rect 56 53 119 54
rect 166 56 278 57
rect 166 54 167 56
rect 169 54 275 56
rect 277 54 278 56
rect 166 53 278 54
rect 341 56 404 57
rect 341 54 342 56
rect 344 54 385 56
rect 387 54 401 56
rect 403 54 404 56
rect 341 53 404 54
rect 488 56 600 57
rect 488 54 489 56
rect 491 54 552 56
rect 554 54 597 56
rect 599 54 600 56
rect 488 53 600 54
rect -699 48 -660 49
rect -699 46 -698 48
rect -696 46 -663 48
rect -661 46 -660 48
rect -699 45 -660 46
rect -648 48 -569 49
rect -648 46 -647 48
rect -645 46 -626 48
rect -624 46 -572 48
rect -570 46 -569 48
rect -648 45 -569 46
rect -363 48 -284 49
rect -363 46 -362 48
rect -360 46 -341 48
rect -339 46 -287 48
rect -285 46 -284 48
rect -363 45 -284 46
rect -78 48 1 49
rect -78 46 -77 48
rect -75 46 -56 48
rect -54 46 -2 48
rect 0 46 1 48
rect -78 45 1 46
rect 207 48 286 49
rect 207 46 208 48
rect 210 46 229 48
rect 231 46 283 48
rect 285 46 286 48
rect 207 45 286 46
rect 454 48 458 49
rect 454 46 455 48
rect 457 46 458 48
rect 454 45 458 46
rect 514 48 518 49
rect 514 46 515 48
rect 517 46 518 48
rect 514 45 518 46
rect 580 48 612 49
rect 580 46 581 48
rect 583 46 609 48
rect 611 46 612 48
rect 580 45 612 46
rect -594 40 -479 41
rect -594 38 -593 40
rect -591 38 -482 40
rect -480 38 -479 40
rect -594 37 -479 38
rect -309 40 -194 41
rect -309 38 -308 40
rect -306 38 -197 40
rect -195 38 -194 40
rect -309 37 -194 38
rect -24 40 91 41
rect -24 38 -23 40
rect -21 38 88 40
rect 90 38 91 40
rect -24 37 91 38
rect 156 40 205 41
rect 156 38 157 40
rect 159 38 202 40
rect 204 38 205 40
rect 156 37 205 38
rect 261 40 376 41
rect 261 38 262 40
rect 264 38 373 40
rect 375 38 376 40
rect 261 37 376 38
rect 538 40 620 41
rect 538 38 539 40
rect 541 38 617 40
rect 619 38 620 40
rect 538 37 620 38
rect 680 33 708 34
rect -664 32 -443 33
rect -664 30 -663 32
rect -661 30 -446 32
rect -444 30 -443 32
rect -664 29 -443 30
rect -379 32 -158 33
rect -379 30 -378 32
rect -376 30 -161 32
rect -159 30 -158 32
rect -379 29 -158 30
rect -94 32 127 33
rect -94 30 -93 32
rect -91 30 124 32
rect 126 30 127 32
rect -94 29 127 30
rect 191 32 412 33
rect 191 30 192 32
rect 194 30 409 32
rect 411 30 412 32
rect 191 29 412 30
rect 478 32 628 33
rect 478 30 479 32
rect 481 30 625 32
rect 627 30 628 32
rect 680 31 681 33
rect 683 31 705 33
rect 707 31 708 33
rect 680 30 708 31
rect 478 29 628 30
rect -618 24 -434 25
rect -618 22 -617 24
rect -615 22 -563 24
rect -561 22 -437 24
rect -435 22 -434 24
rect -618 21 -434 22
rect -333 24 -149 25
rect -333 22 -332 24
rect -330 22 -278 24
rect -276 22 -152 24
rect -150 22 -149 24
rect -333 21 -149 22
rect -48 24 136 25
rect -48 22 -47 24
rect -45 22 7 24
rect 9 22 133 24
rect 135 22 136 24
rect -48 21 136 22
rect 237 24 421 25
rect 237 22 238 24
rect 240 22 292 24
rect 294 22 418 24
rect 420 22 421 24
rect 237 21 421 22
rect 441 24 724 25
rect 441 22 442 24
rect 444 22 721 24
rect 723 22 724 24
rect 441 21 724 22
rect -618 16 458 17
rect -618 14 -617 16
rect -615 14 -332 16
rect -330 14 -47 16
rect -45 14 238 16
rect 240 14 455 16
rect 457 14 458 16
rect -618 13 458 14
rect -664 8 195 9
rect -664 6 -663 8
rect -661 6 -378 8
rect -376 6 -93 8
rect -91 6 192 8
rect 194 6 195 8
rect -664 5 195 6
rect 201 8 684 9
rect 201 6 202 8
rect 204 6 681 8
rect 683 6 684 8
rect 201 5 684 6
rect -414 0 149 1
rect -414 -2 -413 0
rect -411 -2 146 0
rect 148 -2 149 0
rect -414 -3 149 -2
rect 166 0 644 1
rect 166 -2 167 0
rect 169 -2 641 0
rect 643 -2 644 0
rect 166 -3 644 -2
rect -707 -8 -400 -7
rect -707 -10 -706 -8
rect -704 -10 -403 -8
rect -401 -10 -400 -8
rect -707 -11 -400 -10
rect -129 -8 140 -7
rect -129 -10 -128 -8
rect -126 -10 137 -8
rect 139 -10 140 -8
rect -129 -11 140 -10
rect 145 -8 473 -7
rect 145 -10 146 -8
rect 148 -10 470 -8
rect 472 -10 473 -8
rect 145 -11 473 -10
rect -119 -16 652 -15
rect -119 -18 -118 -16
rect -116 -18 649 -16
rect 651 -18 652 -16
rect -119 -19 652 -18
rect -715 -24 -685 -23
rect -715 -26 -714 -24
rect -712 -26 -688 -24
rect -686 -26 -685 -24
rect -715 -27 -685 -26
rect 136 -24 555 -23
rect 136 -26 137 -24
rect 139 -26 552 -24
rect 554 -26 555 -24
rect 136 -27 555 -26
rect -715 -40 -685 -39
rect -715 -42 -714 -40
rect -712 -42 -688 -40
rect -686 -42 -685 -40
rect -715 -43 -685 -42
rect 156 -40 700 -39
rect 156 -42 157 -40
rect 159 -42 697 -40
rect 699 -42 700 -40
rect 156 -43 700 -42
rect -119 -48 652 -47
rect -119 -50 -118 -48
rect -116 -50 649 -48
rect 651 -50 652 -48
rect -119 -51 652 -50
rect -707 -56 -400 -55
rect -707 -58 -706 -56
rect -704 -58 -403 -56
rect -401 -58 -400 -56
rect -707 -59 -400 -58
rect -129 -56 144 -55
rect -129 -58 -128 -56
rect -126 -58 141 -56
rect 143 -58 144 -56
rect -129 -59 144 -58
rect 148 -56 463 -55
rect 148 -58 149 -56
rect 151 -58 460 -56
rect 462 -58 463 -56
rect 148 -59 463 -58
rect -414 -64 152 -63
rect -414 -66 -413 -64
rect -411 -66 149 -64
rect 151 -66 152 -64
rect -414 -67 152 -66
rect 166 -64 644 -63
rect 166 -66 167 -64
rect 169 -66 641 -64
rect 643 -66 644 -64
rect 166 -67 644 -66
rect -664 -72 195 -71
rect -664 -74 -663 -72
rect -661 -74 -378 -72
rect -376 -74 -93 -72
rect -91 -74 192 -72
rect 194 -74 195 -72
rect -664 -75 195 -74
rect 229 -72 565 -71
rect 229 -74 230 -72
rect 232 -74 562 -72
rect 564 -74 565 -72
rect 229 -75 565 -74
rect -618 -80 518 -79
rect -618 -82 -617 -80
rect -615 -82 -332 -80
rect -330 -82 -47 -80
rect -45 -82 238 -80
rect 240 -82 515 -80
rect 517 -82 518 -80
rect -618 -83 518 -82
rect -618 -88 -434 -87
rect -618 -90 -617 -88
rect -615 -90 -563 -88
rect -561 -90 -437 -88
rect -435 -90 -434 -88
rect -618 -91 -434 -90
rect -333 -88 -149 -87
rect -333 -90 -332 -88
rect -330 -90 -278 -88
rect -276 -90 -152 -88
rect -150 -90 -149 -88
rect -333 -91 -149 -90
rect -48 -88 136 -87
rect -48 -90 -47 -88
rect -45 -90 7 -88
rect 9 -90 133 -88
rect 135 -90 136 -88
rect -48 -91 136 -90
rect 140 -88 233 -87
rect 140 -90 141 -88
rect 143 -90 230 -88
rect 232 -90 233 -88
rect 140 -91 233 -90
rect 237 -88 421 -87
rect 237 -90 238 -88
rect 240 -90 292 -88
rect 294 -90 418 -88
rect 420 -90 421 -88
rect 237 -91 421 -90
rect 441 -88 716 -87
rect 441 -90 442 -88
rect 444 -90 713 -88
rect 715 -90 716 -88
rect 441 -91 716 -90
rect -664 -96 -443 -95
rect -664 -98 -663 -96
rect -661 -98 -446 -96
rect -444 -98 -443 -96
rect -664 -99 -443 -98
rect -379 -96 -158 -95
rect -379 -98 -378 -96
rect -376 -98 -161 -96
rect -159 -98 -158 -96
rect -379 -99 -158 -98
rect -94 -96 127 -95
rect -94 -98 -93 -96
rect -91 -98 124 -96
rect 126 -98 127 -96
rect -94 -99 127 -98
rect 191 -96 412 -95
rect 191 -98 192 -96
rect 194 -98 409 -96
rect 411 -98 412 -96
rect 191 -99 412 -98
rect 680 -96 692 -95
rect 680 -98 681 -96
rect 683 -98 689 -96
rect 691 -98 692 -96
rect 680 -99 692 -98
rect -594 -104 -479 -103
rect -594 -106 -593 -104
rect -591 -106 -482 -104
rect -480 -106 -479 -104
rect -594 -107 -479 -106
rect -309 -104 -194 -103
rect -309 -106 -308 -104
rect -306 -106 -197 -104
rect -195 -106 -194 -104
rect -309 -107 -194 -106
rect -24 -104 91 -103
rect -24 -106 -23 -104
rect -21 -106 88 -104
rect 90 -106 91 -104
rect -24 -107 91 -106
rect 261 -104 376 -103
rect 261 -106 262 -104
rect 264 -106 373 -104
rect 375 -106 376 -104
rect 261 -107 376 -106
rect 590 -104 668 -103
rect 590 -106 591 -104
rect 593 -106 665 -104
rect 667 -106 668 -104
rect 590 -107 668 -106
rect 672 -104 684 -103
rect 672 -106 673 -104
rect 675 -106 681 -104
rect 683 -106 684 -104
rect 672 -107 684 -106
rect -699 -112 -660 -111
rect -699 -114 -698 -112
rect -696 -114 -663 -112
rect -661 -114 -660 -112
rect -699 -115 -660 -114
rect -648 -112 -569 -111
rect -648 -114 -647 -112
rect -645 -114 -626 -112
rect -624 -114 -572 -112
rect -570 -114 -569 -112
rect -648 -115 -569 -114
rect -363 -112 -284 -111
rect -363 -114 -362 -112
rect -360 -114 -341 -112
rect -339 -114 -287 -112
rect -285 -114 -284 -112
rect -363 -115 -284 -114
rect -78 -112 1 -111
rect -78 -114 -77 -112
rect -75 -114 -56 -112
rect -54 -114 -2 -112
rect 0 -114 1 -112
rect -78 -115 1 -114
rect 207 -112 286 -111
rect 207 -114 208 -112
rect 210 -114 229 -112
rect 231 -114 283 -112
rect 285 -114 286 -112
rect 207 -115 286 -114
rect 579 -112 676 -111
rect 579 -114 580 -112
rect 582 -114 673 -112
rect 675 -114 676 -112
rect 579 -115 676 -114
rect -689 -120 -577 -119
rect -689 -122 -688 -120
rect -686 -122 -580 -120
rect -578 -122 -577 -120
rect -689 -123 -577 -122
rect -514 -120 -451 -119
rect -514 -122 -513 -120
rect -511 -122 -470 -120
rect -468 -122 -454 -120
rect -452 -122 -451 -120
rect -514 -123 -451 -122
rect -404 -120 -292 -119
rect -404 -122 -403 -120
rect -401 -122 -295 -120
rect -293 -122 -292 -120
rect -404 -123 -292 -122
rect -229 -120 -166 -119
rect -229 -122 -228 -120
rect -226 -122 -185 -120
rect -183 -122 -169 -120
rect -167 -122 -166 -120
rect -229 -123 -166 -122
rect -119 -120 -7 -119
rect -119 -122 -118 -120
rect -116 -122 -10 -120
rect -8 -122 -7 -120
rect -119 -123 -7 -122
rect 56 -120 119 -119
rect 56 -122 57 -120
rect 59 -122 100 -120
rect 102 -122 116 -120
rect 118 -122 119 -120
rect 56 -123 119 -122
rect 166 -120 278 -119
rect 166 -122 167 -120
rect 169 -122 275 -120
rect 277 -122 278 -120
rect 166 -123 278 -122
rect 341 -120 404 -119
rect 341 -122 342 -120
rect 344 -122 385 -120
rect 387 -122 401 -120
rect 403 -122 404 -120
rect 341 -123 404 -122
rect 498 -120 668 -119
rect 498 -122 499 -120
rect 501 -122 665 -120
rect 667 -122 668 -120
rect 498 -123 668 -122
rect -674 -128 -631 -127
rect -674 -130 -673 -128
rect -671 -130 -634 -128
rect -632 -130 -631 -128
rect -674 -131 -631 -130
rect -540 -128 -526 -127
rect -540 -130 -539 -128
rect -537 -130 -529 -128
rect -527 -130 -526 -128
rect -540 -131 -526 -130
rect -506 -128 -491 -127
rect -506 -130 -505 -128
rect -503 -130 -494 -128
rect -492 -130 -491 -128
rect -506 -131 -491 -130
rect -483 -128 -479 -127
rect -483 -130 -482 -128
rect -480 -130 -479 -128
rect -483 -131 -479 -130
rect -389 -128 -346 -127
rect -389 -130 -388 -128
rect -386 -130 -349 -128
rect -347 -130 -346 -128
rect -389 -131 -346 -130
rect -255 -128 -241 -127
rect -255 -130 -254 -128
rect -252 -130 -244 -128
rect -242 -130 -241 -128
rect -255 -131 -241 -130
rect -221 -128 -206 -127
rect -221 -130 -220 -128
rect -218 -130 -209 -128
rect -207 -130 -206 -128
rect -221 -131 -206 -130
rect -198 -128 -194 -127
rect -198 -130 -197 -128
rect -195 -130 -194 -128
rect -198 -131 -194 -130
rect -104 -128 -61 -127
rect -104 -130 -103 -128
rect -101 -130 -64 -128
rect -62 -130 -61 -128
rect -104 -131 -61 -130
rect 30 -128 44 -127
rect 30 -130 31 -128
rect 33 -130 41 -128
rect 43 -130 44 -128
rect 30 -131 44 -130
rect 64 -128 79 -127
rect 64 -130 65 -128
rect 67 -130 76 -128
rect 78 -130 79 -128
rect 64 -131 79 -130
rect 87 -128 91 -127
rect 87 -130 88 -128
rect 90 -130 91 -128
rect 87 -131 91 -130
rect 181 -128 224 -127
rect 181 -130 182 -128
rect 184 -130 221 -128
rect 223 -130 224 -128
rect 181 -131 224 -130
rect 315 -128 329 -127
rect 315 -130 316 -128
rect 318 -130 326 -128
rect 328 -130 329 -128
rect 315 -131 329 -130
rect 349 -128 364 -127
rect 349 -130 350 -128
rect 352 -130 361 -128
rect 363 -130 364 -128
rect 349 -131 364 -130
rect 372 -128 376 -127
rect 372 -130 373 -128
rect 375 -130 376 -128
rect 372 -131 376 -130
rect 487 -128 660 -127
rect 487 -130 488 -128
rect 490 -130 657 -128
rect 659 -130 660 -128
rect 487 -131 660 -130
rect -690 -139 744 -136
rect -690 -141 739 -139
rect 741 -141 744 -139
rect -690 -143 -687 -141
rect -685 -143 -675 -141
rect -673 -143 -661 -141
rect -659 -143 -649 -141
rect -647 -143 -605 -141
rect -603 -143 -595 -141
rect -593 -143 -551 -141
rect -549 -143 -541 -141
rect -539 -143 -527 -141
rect -525 -143 -506 -141
rect -504 -143 -492 -141
rect -490 -143 -471 -141
rect -469 -143 -425 -141
rect -423 -143 -415 -141
rect -413 -143 -402 -141
rect -400 -143 -390 -141
rect -388 -143 -376 -141
rect -374 -143 -364 -141
rect -362 -143 -320 -141
rect -318 -143 -310 -141
rect -308 -143 -266 -141
rect -264 -143 -256 -141
rect -254 -143 -242 -141
rect -240 -143 -221 -141
rect -219 -143 -207 -141
rect -205 -143 -186 -141
rect -184 -143 -140 -141
rect -138 -143 -130 -141
rect -128 -143 -117 -141
rect -115 -143 -105 -141
rect -103 -143 -91 -141
rect -89 -143 -79 -141
rect -77 -143 -35 -141
rect -33 -143 -25 -141
rect -23 -143 19 -141
rect 21 -143 29 -141
rect 31 -143 43 -141
rect 45 -143 64 -141
rect 66 -143 78 -141
rect 80 -143 99 -141
rect 101 -143 145 -141
rect 147 -143 155 -141
rect 157 -143 168 -141
rect 170 -143 180 -141
rect 182 -143 194 -141
rect 196 -143 206 -141
rect 208 -143 250 -141
rect 252 -143 260 -141
rect 262 -143 304 -141
rect 306 -143 314 -141
rect 316 -143 328 -141
rect 330 -143 349 -141
rect 351 -143 363 -141
rect 365 -143 384 -141
rect 386 -143 430 -141
rect 432 -143 440 -141
rect 442 -143 461 -141
rect 463 -143 469 -141
rect 471 -143 479 -141
rect 481 -143 501 -141
rect 503 -143 523 -141
rect 525 -143 553 -141
rect 555 -143 561 -141
rect 563 -143 571 -141
rect 573 -143 593 -141
rect 595 -143 615 -141
rect 617 -143 744 -141
rect -690 -144 744 -143
rect -682 -165 -678 -157
rect -674 -158 -670 -149
rect -672 -160 -670 -158
rect -690 -167 -678 -165
rect -690 -169 -688 -167
rect -686 -169 -681 -167
rect -679 -169 -678 -167
rect -690 -171 -678 -169
rect -674 -164 -670 -160
rect -674 -166 -673 -164
rect -671 -166 -670 -164
rect -656 -165 -652 -157
rect -648 -158 -644 -149
rect -646 -160 -644 -158
rect -674 -176 -670 -166
rect -664 -167 -652 -165
rect -664 -169 -663 -167
rect -661 -169 -655 -167
rect -653 -169 -652 -167
rect -664 -171 -652 -169
rect -648 -164 -644 -160
rect -648 -166 -647 -164
rect -645 -166 -644 -164
rect -672 -178 -670 -176
rect -674 -181 -670 -178
rect -648 -176 -644 -166
rect -635 -158 -622 -157
rect -635 -160 -634 -158
rect -632 -160 -622 -158
rect -635 -163 -622 -160
rect -618 -160 -614 -157
rect -618 -162 -617 -160
rect -615 -162 -614 -160
rect -594 -157 -590 -149
rect -592 -159 -590 -157
rect -635 -167 -629 -163
rect -635 -169 -633 -167
rect -631 -169 -629 -167
rect -635 -170 -629 -169
rect -618 -166 -614 -162
rect -618 -167 -605 -166
rect -618 -169 -611 -167
rect -609 -169 -605 -167
rect -618 -170 -605 -169
rect -646 -178 -644 -176
rect -635 -175 -621 -174
rect -635 -177 -626 -175
rect -624 -176 -621 -175
rect -619 -176 -613 -174
rect -624 -177 -613 -176
rect -635 -178 -613 -177
rect -594 -165 -590 -159
rect -594 -167 -593 -165
rect -591 -167 -590 -165
rect -648 -181 -644 -178
rect -682 -183 -670 -181
rect -682 -185 -674 -183
rect -672 -185 -670 -183
rect -682 -187 -670 -185
rect -656 -183 -644 -181
rect -656 -185 -648 -183
rect -646 -185 -644 -183
rect -656 -187 -644 -185
rect -627 -186 -621 -178
rect -594 -178 -590 -167
rect -581 -158 -568 -157
rect -581 -160 -580 -158
rect -578 -160 -568 -158
rect -581 -163 -568 -160
rect -564 -160 -560 -157
rect -564 -162 -563 -160
rect -561 -162 -560 -160
rect -540 -157 -536 -149
rect -519 -150 -502 -149
rect -519 -152 -517 -150
rect -515 -152 -502 -150
rect -519 -153 -502 -152
rect -514 -155 -502 -153
rect -538 -159 -536 -157
rect -581 -167 -575 -163
rect -581 -169 -579 -167
rect -577 -169 -575 -167
rect -581 -170 -575 -169
rect -564 -166 -560 -162
rect -564 -167 -551 -166
rect -564 -169 -557 -167
rect -555 -169 -551 -167
rect -564 -170 -551 -169
rect -581 -175 -567 -174
rect -581 -177 -572 -175
rect -570 -176 -567 -175
rect -565 -176 -559 -174
rect -570 -177 -559 -176
rect -581 -178 -559 -177
rect -540 -165 -536 -159
rect -522 -163 -518 -157
rect -540 -167 -539 -165
rect -537 -167 -536 -165
rect -592 -180 -590 -178
rect -594 -182 -590 -180
rect -603 -185 -590 -182
rect -603 -186 -594 -185
rect -595 -187 -594 -186
rect -592 -187 -590 -185
rect -595 -195 -590 -187
rect -573 -186 -567 -178
rect -540 -178 -536 -167
rect -530 -164 -518 -163
rect -530 -166 -529 -164
rect -527 -166 -523 -164
rect -521 -166 -518 -164
rect -506 -159 -502 -155
rect -484 -150 -467 -149
rect -484 -152 -482 -150
rect -480 -152 -467 -150
rect -484 -153 -467 -152
rect -479 -155 -467 -153
rect -471 -157 -467 -155
rect -506 -161 -505 -159
rect -503 -161 -502 -159
rect -530 -167 -518 -166
rect -514 -167 -510 -165
rect -530 -171 -526 -167
rect -514 -169 -513 -167
rect -511 -169 -510 -167
rect -514 -171 -510 -169
rect -538 -180 -536 -178
rect -522 -172 -510 -171
rect -522 -174 -513 -172
rect -511 -174 -510 -172
rect -522 -175 -510 -174
rect -522 -179 -518 -175
rect -540 -182 -536 -180
rect -549 -185 -536 -182
rect -506 -183 -502 -161
rect -487 -163 -483 -157
rect -495 -164 -483 -163
rect -495 -166 -494 -164
rect -492 -166 -488 -164
rect -486 -166 -483 -164
rect -471 -159 -470 -157
rect -468 -159 -467 -157
rect -495 -167 -483 -166
rect -479 -167 -475 -165
rect -495 -171 -491 -167
rect -479 -169 -478 -167
rect -476 -169 -475 -167
rect -479 -171 -475 -169
rect -487 -172 -475 -171
rect -487 -174 -482 -172
rect -480 -174 -475 -172
rect -487 -175 -475 -174
rect -487 -179 -483 -175
rect -471 -183 -467 -159
rect -455 -158 -442 -157
rect -455 -160 -454 -158
rect -452 -160 -442 -158
rect -455 -163 -442 -160
rect -438 -159 -434 -157
rect -438 -161 -437 -159
rect -435 -161 -434 -159
rect -414 -157 -410 -149
rect -412 -159 -410 -157
rect -414 -161 -410 -159
rect -455 -167 -449 -163
rect -455 -169 -453 -167
rect -451 -169 -449 -167
rect -455 -170 -449 -169
rect -438 -166 -434 -161
rect -438 -167 -425 -166
rect -438 -169 -431 -167
rect -429 -169 -425 -167
rect -438 -170 -425 -169
rect -455 -175 -441 -174
rect -455 -177 -446 -175
rect -444 -176 -441 -175
rect -439 -176 -433 -174
rect -444 -177 -433 -176
rect -455 -178 -433 -177
rect -414 -163 -413 -161
rect -411 -163 -410 -161
rect -549 -186 -540 -185
rect -541 -187 -540 -186
rect -538 -187 -536 -185
rect -541 -195 -536 -187
rect -511 -184 -502 -183
rect -511 -186 -509 -184
rect -507 -186 -502 -184
rect -511 -187 -502 -186
rect -476 -184 -467 -183
rect -476 -186 -474 -184
rect -472 -186 -467 -184
rect -476 -187 -467 -186
rect -511 -191 -505 -187
rect -511 -193 -509 -191
rect -507 -193 -505 -191
rect -511 -194 -505 -193
rect -476 -191 -470 -187
rect -476 -193 -474 -191
rect -472 -193 -470 -191
rect -476 -194 -470 -193
rect -447 -186 -441 -178
rect -414 -178 -410 -163
rect -397 -165 -393 -157
rect -389 -158 -385 -149
rect -387 -160 -385 -158
rect -405 -167 -393 -165
rect -405 -169 -403 -167
rect -401 -169 -396 -167
rect -394 -169 -393 -167
rect -405 -171 -393 -169
rect -389 -164 -385 -160
rect -389 -166 -388 -164
rect -386 -166 -385 -164
rect -371 -165 -367 -157
rect -363 -158 -359 -149
rect -361 -160 -359 -158
rect -412 -180 -410 -178
rect -414 -182 -410 -180
rect -389 -176 -385 -166
rect -379 -167 -367 -165
rect -379 -169 -378 -167
rect -376 -169 -370 -167
rect -368 -169 -367 -167
rect -379 -171 -367 -169
rect -363 -164 -359 -160
rect -363 -166 -362 -164
rect -360 -166 -359 -164
rect -387 -178 -385 -176
rect -389 -181 -385 -178
rect -363 -176 -359 -166
rect -350 -158 -337 -157
rect -350 -160 -349 -158
rect -347 -160 -337 -158
rect -350 -163 -337 -160
rect -333 -160 -329 -157
rect -333 -162 -332 -160
rect -330 -162 -329 -160
rect -309 -157 -305 -149
rect -307 -159 -305 -157
rect -350 -167 -344 -163
rect -350 -169 -348 -167
rect -346 -169 -344 -167
rect -350 -170 -344 -169
rect -333 -166 -329 -162
rect -333 -167 -320 -166
rect -333 -169 -326 -167
rect -324 -169 -320 -167
rect -333 -170 -320 -169
rect -361 -178 -359 -176
rect -350 -175 -336 -174
rect -350 -177 -341 -175
rect -339 -176 -336 -175
rect -334 -176 -328 -174
rect -339 -177 -328 -176
rect -350 -178 -328 -177
rect -309 -165 -305 -159
rect -309 -167 -308 -165
rect -306 -167 -305 -165
rect -363 -181 -359 -178
rect -423 -185 -410 -182
rect -423 -186 -414 -185
rect -415 -187 -414 -186
rect -412 -187 -410 -185
rect -397 -183 -385 -181
rect -397 -185 -389 -183
rect -387 -185 -385 -183
rect -397 -187 -385 -185
rect -371 -183 -359 -181
rect -371 -185 -363 -183
rect -361 -185 -359 -183
rect -371 -187 -359 -185
rect -471 -200 -464 -199
rect -415 -195 -410 -187
rect -342 -186 -336 -178
rect -309 -178 -305 -167
rect -296 -158 -283 -157
rect -296 -160 -295 -158
rect -293 -160 -283 -158
rect -296 -163 -283 -160
rect -279 -160 -275 -157
rect -279 -162 -278 -160
rect -276 -162 -275 -160
rect -255 -157 -251 -149
rect -234 -150 -217 -149
rect -234 -152 -232 -150
rect -230 -152 -217 -150
rect -234 -153 -217 -152
rect -229 -155 -217 -153
rect -253 -159 -251 -157
rect -296 -167 -290 -163
rect -296 -169 -294 -167
rect -292 -169 -290 -167
rect -296 -170 -290 -169
rect -279 -166 -275 -162
rect -279 -167 -266 -166
rect -279 -169 -272 -167
rect -270 -169 -266 -167
rect -279 -170 -266 -169
rect -296 -175 -282 -174
rect -296 -177 -287 -175
rect -285 -176 -282 -175
rect -280 -176 -274 -174
rect -285 -177 -274 -176
rect -296 -178 -274 -177
rect -255 -165 -251 -159
rect -237 -163 -233 -157
rect -255 -167 -254 -165
rect -252 -167 -251 -165
rect -307 -180 -305 -178
rect -309 -182 -305 -180
rect -318 -185 -305 -182
rect -318 -186 -309 -185
rect -310 -187 -309 -186
rect -307 -187 -305 -185
rect -310 -195 -305 -187
rect -288 -186 -282 -178
rect -255 -178 -251 -167
rect -245 -164 -233 -163
rect -245 -166 -244 -164
rect -242 -166 -238 -164
rect -236 -166 -233 -164
rect -221 -159 -217 -155
rect -199 -150 -182 -149
rect -199 -152 -197 -150
rect -195 -152 -182 -150
rect -199 -153 -182 -152
rect -194 -155 -182 -153
rect -186 -157 -182 -155
rect -221 -161 -220 -159
rect -218 -161 -217 -159
rect -245 -167 -233 -166
rect -229 -167 -225 -165
rect -245 -171 -241 -167
rect -229 -169 -228 -167
rect -226 -169 -225 -167
rect -229 -171 -225 -169
rect -253 -180 -251 -178
rect -237 -172 -225 -171
rect -237 -174 -228 -172
rect -226 -174 -225 -172
rect -237 -175 -225 -174
rect -237 -179 -233 -175
rect -255 -182 -251 -180
rect -264 -185 -251 -182
rect -221 -183 -217 -161
rect -202 -163 -198 -157
rect -210 -164 -198 -163
rect -210 -166 -209 -164
rect -207 -166 -203 -164
rect -201 -166 -198 -164
rect -186 -159 -185 -157
rect -183 -159 -182 -157
rect -210 -167 -198 -166
rect -194 -167 -190 -165
rect -210 -171 -206 -167
rect -194 -169 -193 -167
rect -191 -169 -190 -167
rect -194 -171 -190 -169
rect -202 -172 -190 -171
rect -202 -174 -197 -172
rect -195 -174 -190 -172
rect -202 -175 -190 -174
rect -202 -179 -198 -175
rect -186 -183 -182 -159
rect -170 -158 -157 -157
rect -170 -160 -169 -158
rect -167 -160 -157 -158
rect -170 -163 -157 -160
rect -153 -159 -149 -157
rect -153 -161 -152 -159
rect -150 -161 -149 -159
rect -129 -157 -125 -149
rect -127 -159 -125 -157
rect -129 -161 -125 -159
rect -170 -167 -164 -163
rect -170 -169 -168 -167
rect -166 -169 -164 -167
rect -170 -170 -164 -169
rect -153 -166 -149 -161
rect -153 -167 -140 -166
rect -153 -169 -146 -167
rect -144 -169 -140 -167
rect -153 -170 -140 -169
rect -170 -175 -156 -174
rect -170 -177 -161 -175
rect -159 -176 -156 -175
rect -154 -176 -148 -174
rect -159 -177 -148 -176
rect -170 -178 -148 -177
rect -129 -163 -128 -161
rect -126 -163 -125 -161
rect -264 -186 -255 -185
rect -256 -187 -255 -186
rect -253 -187 -251 -185
rect -256 -195 -251 -187
rect -226 -184 -217 -183
rect -226 -186 -224 -184
rect -222 -186 -217 -184
rect -226 -187 -217 -186
rect -191 -184 -182 -183
rect -191 -186 -189 -184
rect -187 -186 -182 -184
rect -191 -187 -182 -186
rect -226 -191 -220 -187
rect -226 -193 -224 -191
rect -222 -193 -220 -191
rect -226 -194 -220 -193
rect -191 -191 -185 -187
rect -191 -193 -189 -191
rect -187 -193 -185 -191
rect -191 -194 -185 -193
rect -162 -186 -156 -178
rect -129 -178 -125 -163
rect -112 -165 -108 -157
rect -104 -158 -100 -149
rect -102 -160 -100 -158
rect -120 -167 -108 -165
rect -120 -169 -118 -167
rect -116 -169 -111 -167
rect -109 -169 -108 -167
rect -120 -171 -108 -169
rect -104 -164 -100 -160
rect -104 -166 -103 -164
rect -101 -166 -100 -164
rect -86 -165 -82 -157
rect -78 -158 -74 -149
rect -76 -160 -74 -158
rect -127 -180 -125 -178
rect -129 -182 -125 -180
rect -104 -176 -100 -166
rect -94 -167 -82 -165
rect -94 -169 -93 -167
rect -91 -169 -85 -167
rect -83 -169 -82 -167
rect -94 -171 -82 -169
rect -78 -164 -74 -160
rect -78 -166 -77 -164
rect -75 -166 -74 -164
rect -102 -178 -100 -176
rect -104 -181 -100 -178
rect -78 -176 -74 -166
rect -65 -158 -52 -157
rect -65 -160 -64 -158
rect -62 -160 -52 -158
rect -65 -163 -52 -160
rect -48 -160 -44 -157
rect -48 -162 -47 -160
rect -45 -162 -44 -160
rect -24 -157 -20 -149
rect -22 -159 -20 -157
rect -65 -167 -59 -163
rect -65 -169 -63 -167
rect -61 -169 -59 -167
rect -65 -170 -59 -169
rect -48 -166 -44 -162
rect -48 -167 -35 -166
rect -48 -169 -41 -167
rect -39 -169 -35 -167
rect -48 -170 -35 -169
rect -76 -178 -74 -176
rect -65 -175 -51 -174
rect -65 -177 -56 -175
rect -54 -176 -51 -175
rect -49 -176 -43 -174
rect -54 -177 -43 -176
rect -65 -178 -43 -177
rect -24 -165 -20 -159
rect -24 -167 -23 -165
rect -21 -167 -20 -165
rect -78 -181 -74 -178
rect -138 -185 -125 -182
rect -138 -186 -129 -185
rect -130 -187 -129 -186
rect -127 -187 -125 -185
rect -112 -183 -100 -181
rect -112 -185 -104 -183
rect -102 -185 -100 -183
rect -112 -187 -100 -185
rect -86 -183 -74 -181
rect -86 -185 -78 -183
rect -76 -185 -74 -183
rect -86 -187 -74 -185
rect -186 -200 -179 -199
rect -130 -195 -125 -187
rect -57 -186 -51 -178
rect -24 -178 -20 -167
rect -11 -158 2 -157
rect -11 -160 -10 -158
rect -8 -160 2 -158
rect -11 -163 2 -160
rect 6 -160 10 -157
rect 6 -162 7 -160
rect 9 -162 10 -160
rect 30 -157 34 -149
rect 51 -150 68 -149
rect 51 -152 53 -150
rect 55 -152 68 -150
rect 51 -153 68 -152
rect 56 -155 68 -153
rect 32 -159 34 -157
rect -11 -167 -5 -163
rect -11 -169 -9 -167
rect -7 -169 -5 -167
rect -11 -170 -5 -169
rect 6 -166 10 -162
rect 6 -167 19 -166
rect 6 -169 13 -167
rect 15 -169 19 -167
rect 6 -170 19 -169
rect -11 -175 3 -174
rect -11 -177 -2 -175
rect 0 -176 3 -175
rect 5 -176 11 -174
rect 0 -177 11 -176
rect -11 -178 11 -177
rect 30 -165 34 -159
rect 48 -163 52 -157
rect 30 -167 31 -165
rect 33 -167 34 -165
rect -22 -180 -20 -178
rect -24 -182 -20 -180
rect -33 -185 -20 -182
rect -33 -186 -24 -185
rect -25 -187 -24 -186
rect -22 -187 -20 -185
rect -25 -195 -20 -187
rect -3 -186 3 -178
rect 30 -178 34 -167
rect 40 -164 52 -163
rect 40 -166 41 -164
rect 43 -166 47 -164
rect 49 -166 52 -164
rect 64 -159 68 -155
rect 86 -150 103 -149
rect 86 -152 88 -150
rect 90 -152 103 -150
rect 86 -153 103 -152
rect 91 -155 103 -153
rect 99 -157 103 -155
rect 64 -161 65 -159
rect 67 -161 68 -159
rect 40 -167 52 -166
rect 56 -167 60 -165
rect 40 -171 44 -167
rect 56 -169 57 -167
rect 59 -169 60 -167
rect 56 -171 60 -169
rect 32 -180 34 -178
rect 48 -172 60 -171
rect 48 -174 57 -172
rect 59 -174 60 -172
rect 48 -175 60 -174
rect 48 -179 52 -175
rect 30 -182 34 -180
rect 21 -185 34 -182
rect 64 -183 68 -161
rect 83 -163 87 -157
rect 75 -164 87 -163
rect 75 -166 76 -164
rect 78 -166 82 -164
rect 84 -166 87 -164
rect 99 -159 100 -157
rect 102 -159 103 -157
rect 75 -167 87 -166
rect 91 -167 95 -165
rect 75 -171 79 -167
rect 91 -169 92 -167
rect 94 -169 95 -167
rect 91 -171 95 -169
rect 83 -172 95 -171
rect 83 -174 88 -172
rect 90 -174 95 -172
rect 83 -175 95 -174
rect 83 -179 87 -175
rect 99 -183 103 -159
rect 115 -158 128 -157
rect 115 -160 116 -158
rect 118 -160 128 -158
rect 115 -163 128 -160
rect 132 -159 136 -157
rect 132 -161 133 -159
rect 135 -161 136 -159
rect 156 -157 160 -149
rect 158 -159 160 -157
rect 156 -161 160 -159
rect 115 -167 121 -163
rect 115 -169 117 -167
rect 119 -169 121 -167
rect 115 -170 121 -169
rect 132 -166 136 -161
rect 132 -167 145 -166
rect 132 -169 139 -167
rect 141 -169 145 -167
rect 132 -170 145 -169
rect 115 -175 129 -174
rect 115 -177 124 -175
rect 126 -176 129 -175
rect 131 -176 137 -174
rect 126 -177 137 -176
rect 115 -178 137 -177
rect 156 -163 157 -161
rect 159 -163 160 -161
rect 21 -186 30 -185
rect 29 -187 30 -186
rect 32 -187 34 -185
rect 29 -195 34 -187
rect 59 -184 68 -183
rect 59 -186 61 -184
rect 63 -186 68 -184
rect 59 -187 68 -186
rect 94 -184 103 -183
rect 94 -186 96 -184
rect 98 -186 103 -184
rect 94 -187 103 -186
rect 59 -191 65 -187
rect 59 -193 61 -191
rect 63 -193 65 -191
rect 59 -194 65 -193
rect 94 -191 100 -187
rect 94 -193 96 -191
rect 98 -193 100 -191
rect 94 -194 100 -193
rect 123 -186 129 -178
rect 156 -178 160 -163
rect 173 -165 177 -157
rect 181 -158 185 -149
rect 183 -160 185 -158
rect 165 -167 177 -165
rect 165 -169 167 -167
rect 169 -169 174 -167
rect 176 -169 177 -167
rect 165 -171 177 -169
rect 181 -164 185 -160
rect 181 -166 182 -164
rect 184 -166 185 -164
rect 199 -165 203 -157
rect 207 -158 211 -149
rect 209 -160 211 -158
rect 158 -180 160 -178
rect 156 -182 160 -180
rect 181 -176 185 -166
rect 191 -167 203 -165
rect 191 -169 192 -167
rect 194 -169 200 -167
rect 202 -169 203 -167
rect 191 -171 203 -169
rect 207 -164 211 -160
rect 207 -166 208 -164
rect 210 -166 211 -164
rect 183 -178 185 -176
rect 181 -181 185 -178
rect 207 -176 211 -166
rect 220 -158 233 -157
rect 220 -160 221 -158
rect 223 -160 233 -158
rect 220 -163 233 -160
rect 237 -160 241 -157
rect 237 -162 238 -160
rect 240 -162 241 -160
rect 261 -157 265 -149
rect 263 -159 265 -157
rect 220 -167 226 -163
rect 220 -169 222 -167
rect 224 -169 226 -167
rect 220 -170 226 -169
rect 237 -166 241 -162
rect 237 -167 250 -166
rect 237 -169 244 -167
rect 246 -169 250 -167
rect 237 -170 250 -169
rect 209 -178 211 -176
rect 220 -175 234 -174
rect 220 -177 229 -175
rect 231 -176 234 -175
rect 236 -176 242 -174
rect 231 -177 242 -176
rect 220 -178 242 -177
rect 261 -165 265 -159
rect 261 -167 262 -165
rect 264 -167 265 -165
rect 207 -181 211 -178
rect 147 -185 160 -182
rect 147 -186 156 -185
rect 155 -187 156 -186
rect 158 -187 160 -185
rect 173 -183 185 -181
rect 173 -185 181 -183
rect 183 -185 185 -183
rect 173 -187 185 -185
rect 199 -183 211 -181
rect 199 -185 207 -183
rect 209 -185 211 -183
rect 199 -187 211 -185
rect 99 -200 106 -199
rect 155 -195 160 -187
rect 228 -186 234 -178
rect 261 -178 265 -167
rect 274 -158 287 -157
rect 274 -160 275 -158
rect 277 -160 287 -158
rect 274 -163 287 -160
rect 291 -160 295 -157
rect 291 -162 292 -160
rect 294 -162 295 -160
rect 315 -157 319 -149
rect 336 -150 353 -149
rect 336 -152 338 -150
rect 340 -152 353 -150
rect 336 -153 353 -152
rect 341 -155 353 -153
rect 317 -159 319 -157
rect 274 -167 280 -163
rect 274 -169 276 -167
rect 278 -169 280 -167
rect 274 -170 280 -169
rect 291 -166 295 -162
rect 291 -167 304 -166
rect 291 -169 298 -167
rect 300 -169 304 -167
rect 291 -170 304 -169
rect 274 -175 288 -174
rect 274 -177 283 -175
rect 285 -176 288 -175
rect 290 -176 296 -174
rect 285 -177 296 -176
rect 274 -178 296 -177
rect 315 -165 319 -159
rect 333 -163 337 -157
rect 315 -167 316 -165
rect 318 -167 319 -165
rect 263 -180 265 -178
rect 261 -182 265 -180
rect 252 -185 265 -182
rect 252 -186 261 -185
rect 260 -187 261 -186
rect 263 -187 265 -185
rect 260 -195 265 -187
rect 282 -186 288 -178
rect 315 -178 319 -167
rect 325 -164 337 -163
rect 325 -166 326 -164
rect 328 -166 332 -164
rect 334 -166 337 -164
rect 349 -159 353 -155
rect 371 -150 388 -149
rect 371 -152 373 -150
rect 375 -152 388 -150
rect 371 -153 388 -152
rect 376 -155 388 -153
rect 384 -157 388 -155
rect 349 -161 350 -159
rect 352 -161 353 -159
rect 325 -167 337 -166
rect 341 -167 345 -165
rect 325 -171 329 -167
rect 341 -169 342 -167
rect 344 -169 345 -167
rect 341 -171 345 -169
rect 317 -180 319 -178
rect 333 -172 345 -171
rect 333 -174 342 -172
rect 344 -174 345 -172
rect 333 -175 345 -174
rect 333 -179 337 -175
rect 315 -182 319 -180
rect 306 -185 319 -182
rect 349 -183 353 -161
rect 368 -163 372 -157
rect 360 -164 372 -163
rect 360 -166 361 -164
rect 363 -166 367 -164
rect 369 -166 372 -164
rect 384 -159 385 -157
rect 387 -159 388 -157
rect 360 -167 372 -166
rect 376 -167 380 -165
rect 360 -171 364 -167
rect 376 -169 377 -167
rect 379 -169 380 -167
rect 376 -171 380 -169
rect 368 -172 380 -171
rect 368 -174 373 -172
rect 375 -174 380 -172
rect 368 -175 380 -174
rect 368 -179 372 -175
rect 384 -183 388 -159
rect 400 -158 413 -157
rect 400 -160 401 -158
rect 403 -160 413 -158
rect 400 -163 413 -160
rect 417 -159 421 -157
rect 417 -161 418 -159
rect 420 -161 421 -159
rect 441 -157 445 -149
rect 443 -159 445 -157
rect 478 -158 482 -149
rect 441 -161 445 -159
rect 400 -167 406 -163
rect 400 -169 402 -167
rect 404 -169 406 -167
rect 400 -170 406 -169
rect 417 -166 421 -161
rect 417 -167 430 -166
rect 417 -169 424 -167
rect 426 -169 430 -167
rect 417 -170 430 -169
rect 400 -175 414 -174
rect 400 -177 409 -175
rect 411 -176 414 -175
rect 416 -176 422 -174
rect 411 -177 422 -176
rect 400 -178 422 -177
rect 441 -163 442 -161
rect 444 -163 445 -161
rect 475 -159 497 -158
rect 475 -161 477 -159
rect 479 -161 488 -159
rect 490 -161 493 -159
rect 495 -161 497 -159
rect 475 -162 497 -161
rect 306 -186 315 -185
rect 314 -187 315 -186
rect 317 -187 319 -185
rect 314 -195 319 -187
rect 344 -184 353 -183
rect 344 -186 346 -184
rect 348 -186 353 -184
rect 344 -187 353 -186
rect 379 -184 388 -183
rect 379 -186 381 -184
rect 383 -186 388 -184
rect 379 -187 388 -186
rect 344 -191 350 -187
rect 344 -193 346 -191
rect 348 -193 350 -191
rect 344 -194 350 -193
rect 379 -191 385 -187
rect 379 -193 381 -191
rect 383 -193 385 -191
rect 379 -194 385 -193
rect 408 -186 414 -178
rect 441 -178 445 -163
rect 502 -163 506 -157
rect 502 -165 503 -163
rect 505 -165 506 -163
rect 524 -150 538 -149
rect 524 -152 534 -150
rect 536 -152 538 -150
rect 524 -154 538 -152
rect 502 -166 506 -165
rect 469 -169 506 -166
rect 469 -171 471 -169
rect 473 -170 506 -169
rect 473 -171 475 -170
rect 469 -174 475 -171
rect 510 -174 514 -165
rect 443 -180 445 -178
rect 441 -182 445 -180
rect 432 -185 445 -182
rect 432 -186 441 -185
rect 440 -187 441 -186
rect 443 -187 445 -185
rect 459 -175 465 -174
rect 459 -177 461 -175
rect 463 -177 465 -175
rect 459 -179 465 -177
rect 469 -176 470 -174
rect 472 -176 475 -174
rect 469 -178 475 -176
rect 485 -175 514 -174
rect 485 -177 487 -175
rect 489 -177 499 -175
rect 501 -177 514 -175
rect 485 -178 514 -177
rect 459 -181 460 -179
rect 462 -181 465 -179
rect 459 -182 465 -181
rect 518 -173 522 -171
rect 520 -175 522 -173
rect 518 -182 522 -175
rect 459 -186 522 -182
rect 384 -200 391 -199
rect 440 -195 445 -187
rect 478 -195 482 -186
rect 534 -162 538 -154
rect 570 -158 574 -149
rect 567 -159 589 -158
rect 567 -161 569 -159
rect 571 -161 580 -159
rect 582 -161 585 -159
rect 587 -161 589 -159
rect 567 -162 589 -161
rect 534 -164 535 -162
rect 537 -164 538 -162
rect 534 -176 538 -164
rect 594 -163 598 -157
rect 594 -165 595 -163
rect 597 -165 598 -163
rect 616 -150 630 -149
rect 616 -152 626 -150
rect 628 -152 630 -150
rect 616 -154 630 -152
rect 656 -150 708 -149
rect 656 -152 657 -150
rect 659 -152 705 -150
rect 707 -152 708 -150
rect 656 -153 708 -152
rect 594 -166 598 -165
rect 561 -169 598 -166
rect 561 -171 563 -169
rect 565 -170 598 -169
rect 565 -171 567 -170
rect 561 -174 567 -171
rect 602 -174 606 -165
rect 536 -178 538 -176
rect 534 -183 538 -178
rect 536 -185 538 -183
rect 534 -195 538 -185
rect 551 -175 557 -174
rect 551 -177 553 -175
rect 555 -177 557 -175
rect 551 -180 557 -177
rect 561 -176 562 -174
rect 564 -176 567 -174
rect 561 -178 567 -176
rect 577 -175 606 -174
rect 577 -177 579 -175
rect 581 -177 591 -175
rect 593 -177 606 -175
rect 577 -178 606 -177
rect 551 -182 552 -180
rect 554 -182 557 -180
rect 610 -173 614 -171
rect 612 -175 614 -173
rect 610 -182 614 -175
rect 551 -186 614 -182
rect 570 -195 574 -186
rect 626 -176 630 -154
rect 704 -158 716 -157
rect 704 -160 705 -158
rect 707 -160 713 -158
rect 715 -160 716 -158
rect 704 -161 716 -160
rect 712 -166 724 -165
rect 712 -168 713 -166
rect 715 -168 721 -166
rect 723 -168 724 -166
rect 712 -169 724 -168
rect 628 -178 630 -176
rect 626 -183 630 -178
rect 628 -185 630 -183
rect 626 -195 630 -185
rect -738 -201 634 -200
rect -738 -203 -687 -201
rect -685 -203 -675 -201
rect -673 -203 -661 -201
rect -659 -203 -649 -201
rect -647 -203 -639 -201
rect -637 -203 -625 -201
rect -623 -203 -585 -201
rect -583 -203 -571 -201
rect -569 -203 -459 -201
rect -457 -203 -445 -201
rect -443 -203 -402 -201
rect -400 -203 -390 -201
rect -388 -203 -376 -201
rect -374 -203 -364 -201
rect -362 -203 -354 -201
rect -352 -203 -340 -201
rect -338 -203 -300 -201
rect -298 -203 -286 -201
rect -284 -203 -174 -201
rect -172 -203 -160 -201
rect -158 -203 -117 -201
rect -115 -203 -105 -201
rect -103 -203 -91 -201
rect -89 -203 -79 -201
rect -77 -203 -69 -201
rect -67 -203 -55 -201
rect -53 -203 -15 -201
rect -13 -203 -1 -201
rect 1 -203 111 -201
rect 113 -203 125 -201
rect 127 -203 168 -201
rect 170 -203 180 -201
rect 182 -203 194 -201
rect 196 -203 206 -201
rect 208 -203 216 -201
rect 218 -203 230 -201
rect 232 -203 270 -201
rect 272 -203 284 -201
rect 286 -203 396 -201
rect 398 -203 410 -201
rect 412 -203 533 -201
rect 535 -203 625 -201
rect 627 -203 634 -201
rect -738 -207 634 -203
rect -738 -209 -733 -207
rect -731 -209 634 -207
rect -738 -213 634 -209
rect -738 -215 -687 -213
rect -685 -215 -675 -213
rect -673 -215 -661 -213
rect -659 -215 -649 -213
rect -647 -215 -639 -213
rect -637 -215 -625 -213
rect -623 -215 -585 -213
rect -583 -215 -571 -213
rect -569 -215 -459 -213
rect -457 -215 -445 -213
rect -443 -215 -402 -213
rect -400 -215 -390 -213
rect -388 -215 -376 -213
rect -374 -215 -364 -213
rect -362 -215 -354 -213
rect -352 -215 -340 -213
rect -338 -215 -300 -213
rect -298 -215 -286 -213
rect -284 -215 -174 -213
rect -172 -215 -160 -213
rect -158 -215 -117 -213
rect -115 -215 -105 -213
rect -103 -215 -91 -213
rect -89 -215 -79 -213
rect -77 -215 -69 -213
rect -67 -215 -55 -213
rect -53 -215 -15 -213
rect -13 -215 -1 -213
rect 1 -215 111 -213
rect 113 -215 125 -213
rect 127 -215 168 -213
rect 170 -215 180 -213
rect 182 -215 194 -213
rect 196 -215 206 -213
rect 208 -215 216 -213
rect 218 -215 230 -213
rect 232 -215 270 -213
rect 272 -215 284 -213
rect 286 -215 396 -213
rect 398 -215 410 -213
rect 412 -215 533 -213
rect 535 -215 625 -213
rect 627 -215 634 -213
rect -738 -216 634 -215
rect -682 -231 -670 -229
rect -682 -233 -674 -231
rect -672 -233 -670 -231
rect -682 -235 -670 -233
rect -656 -231 -644 -229
rect -656 -233 -648 -231
rect -646 -233 -644 -231
rect -656 -235 -644 -233
rect -674 -238 -670 -235
rect -672 -240 -670 -238
rect -690 -247 -678 -245
rect -690 -249 -688 -247
rect -686 -249 -681 -247
rect -679 -249 -678 -247
rect -690 -251 -678 -249
rect -682 -259 -678 -251
rect -674 -250 -670 -240
rect -648 -238 -644 -235
rect -627 -238 -621 -230
rect -595 -229 -590 -221
rect -595 -230 -594 -229
rect -603 -231 -594 -230
rect -592 -231 -590 -229
rect -603 -234 -590 -231
rect -646 -240 -644 -238
rect -674 -252 -673 -250
rect -671 -252 -670 -250
rect -664 -247 -652 -245
rect -664 -249 -663 -247
rect -661 -249 -655 -247
rect -653 -249 -652 -247
rect -664 -251 -652 -249
rect -674 -256 -670 -252
rect -672 -258 -670 -256
rect -674 -267 -670 -258
rect -656 -259 -652 -251
rect -648 -250 -644 -240
rect -635 -239 -613 -238
rect -635 -241 -626 -239
rect -624 -240 -613 -239
rect -624 -241 -621 -240
rect -635 -242 -621 -241
rect -619 -242 -613 -240
rect -594 -236 -590 -234
rect -592 -238 -590 -236
rect -573 -238 -567 -230
rect -541 -229 -536 -221
rect -471 -217 -464 -216
rect -511 -223 -505 -222
rect -511 -225 -509 -223
rect -507 -225 -505 -223
rect -541 -230 -540 -229
rect -549 -231 -540 -230
rect -538 -231 -536 -229
rect -549 -234 -536 -231
rect -511 -229 -505 -225
rect -476 -223 -470 -222
rect -476 -225 -474 -223
rect -472 -225 -470 -223
rect -476 -229 -470 -225
rect -511 -230 -502 -229
rect -511 -232 -509 -230
rect -507 -232 -502 -230
rect -511 -233 -502 -232
rect -476 -230 -467 -229
rect -476 -232 -474 -230
rect -472 -232 -467 -230
rect -476 -233 -467 -232
rect -648 -252 -647 -250
rect -645 -252 -644 -250
rect -648 -256 -644 -252
rect -646 -258 -644 -256
rect -648 -267 -644 -258
rect -635 -247 -629 -246
rect -635 -249 -633 -247
rect -631 -249 -629 -247
rect -635 -253 -629 -249
rect -618 -247 -605 -246
rect -618 -249 -611 -247
rect -609 -249 -605 -247
rect -618 -250 -605 -249
rect -635 -256 -622 -253
rect -635 -258 -634 -256
rect -632 -258 -622 -256
rect -635 -259 -622 -258
rect -618 -254 -614 -250
rect -618 -256 -617 -254
rect -615 -256 -614 -254
rect -594 -249 -590 -238
rect -581 -239 -559 -238
rect -581 -241 -572 -239
rect -570 -240 -559 -239
rect -570 -241 -567 -240
rect -581 -242 -567 -241
rect -565 -242 -559 -240
rect -540 -236 -536 -234
rect -538 -238 -536 -236
rect -594 -251 -593 -249
rect -591 -251 -590 -249
rect -618 -259 -614 -256
rect -594 -257 -590 -251
rect -592 -259 -590 -257
rect -581 -247 -575 -246
rect -581 -249 -579 -247
rect -577 -249 -575 -247
rect -581 -253 -575 -249
rect -564 -247 -551 -246
rect -564 -249 -557 -247
rect -555 -249 -551 -247
rect -564 -250 -551 -249
rect -581 -256 -568 -253
rect -581 -258 -580 -256
rect -578 -258 -568 -256
rect -581 -259 -568 -258
rect -564 -254 -560 -250
rect -564 -256 -563 -254
rect -561 -256 -560 -254
rect -540 -249 -536 -238
rect -522 -241 -518 -237
rect -522 -242 -510 -241
rect -522 -244 -513 -242
rect -511 -244 -510 -242
rect -522 -245 -510 -244
rect -540 -251 -539 -249
rect -537 -251 -536 -249
rect -564 -259 -560 -256
rect -594 -267 -590 -259
rect -540 -257 -536 -251
rect -530 -249 -526 -245
rect -514 -247 -510 -245
rect -514 -249 -513 -247
rect -511 -249 -510 -247
rect -530 -250 -518 -249
rect -530 -252 -529 -250
rect -527 -252 -523 -250
rect -521 -252 -518 -250
rect -514 -251 -510 -249
rect -530 -253 -518 -252
rect -538 -259 -536 -257
rect -522 -259 -518 -253
rect -506 -255 -502 -233
rect -487 -241 -483 -237
rect -487 -242 -475 -241
rect -487 -244 -482 -242
rect -480 -244 -475 -242
rect -487 -245 -475 -244
rect -495 -249 -491 -245
rect -479 -247 -475 -245
rect -479 -249 -478 -247
rect -476 -249 -475 -247
rect -495 -250 -483 -249
rect -495 -252 -494 -250
rect -492 -252 -488 -250
rect -486 -252 -483 -250
rect -479 -251 -475 -249
rect -495 -253 -483 -252
rect -506 -257 -505 -255
rect -503 -257 -502 -255
rect -540 -267 -536 -259
rect -506 -261 -502 -257
rect -487 -259 -483 -253
rect -471 -257 -467 -233
rect -447 -238 -441 -230
rect -415 -229 -410 -221
rect -415 -230 -414 -229
rect -423 -231 -414 -230
rect -412 -231 -410 -229
rect -423 -234 -410 -231
rect -455 -239 -433 -238
rect -455 -241 -446 -239
rect -444 -240 -433 -239
rect -444 -241 -441 -240
rect -455 -242 -441 -241
rect -439 -242 -433 -240
rect -414 -236 -410 -234
rect -397 -231 -385 -229
rect -397 -233 -389 -231
rect -387 -233 -385 -231
rect -397 -235 -385 -233
rect -371 -231 -359 -229
rect -371 -233 -363 -231
rect -361 -233 -359 -231
rect -371 -235 -359 -233
rect -412 -238 -410 -236
rect -471 -259 -470 -257
rect -468 -259 -467 -257
rect -455 -247 -449 -246
rect -455 -249 -453 -247
rect -451 -249 -449 -247
rect -455 -253 -449 -249
rect -438 -247 -425 -246
rect -438 -249 -431 -247
rect -429 -249 -425 -247
rect -438 -250 -425 -249
rect -455 -256 -442 -253
rect -455 -258 -454 -256
rect -452 -258 -442 -256
rect -455 -259 -442 -258
rect -438 -255 -434 -250
rect -414 -253 -410 -238
rect -389 -238 -385 -235
rect -387 -240 -385 -238
rect -405 -247 -393 -245
rect -405 -249 -403 -247
rect -401 -249 -396 -247
rect -394 -249 -393 -247
rect -405 -251 -393 -249
rect -414 -255 -413 -253
rect -411 -255 -410 -253
rect -438 -257 -437 -255
rect -435 -257 -434 -255
rect -438 -259 -434 -257
rect -514 -263 -502 -261
rect -519 -264 -502 -263
rect -519 -266 -517 -264
rect -515 -266 -502 -264
rect -519 -267 -502 -266
rect -471 -261 -467 -259
rect -479 -263 -467 -261
rect -414 -257 -410 -255
rect -412 -259 -410 -257
rect -484 -264 -467 -263
rect -484 -266 -482 -264
rect -480 -266 -467 -264
rect -484 -267 -467 -266
rect -414 -267 -410 -259
rect -397 -259 -393 -251
rect -389 -250 -385 -240
rect -363 -238 -359 -235
rect -342 -238 -336 -230
rect -310 -229 -305 -221
rect -310 -230 -309 -229
rect -318 -231 -309 -230
rect -307 -231 -305 -229
rect -318 -234 -305 -231
rect -361 -240 -359 -238
rect -389 -252 -388 -250
rect -386 -252 -385 -250
rect -379 -247 -367 -245
rect -379 -249 -378 -247
rect -376 -249 -370 -247
rect -368 -249 -367 -247
rect -379 -251 -367 -249
rect -389 -256 -385 -252
rect -387 -258 -385 -256
rect -389 -267 -385 -258
rect -371 -259 -367 -251
rect -363 -250 -359 -240
rect -350 -239 -328 -238
rect -350 -241 -341 -239
rect -339 -240 -328 -239
rect -339 -241 -336 -240
rect -350 -242 -336 -241
rect -334 -242 -328 -240
rect -309 -236 -305 -234
rect -307 -238 -305 -236
rect -288 -238 -282 -230
rect -256 -229 -251 -221
rect -186 -217 -179 -216
rect -226 -223 -220 -222
rect -226 -225 -224 -223
rect -222 -225 -220 -223
rect -256 -230 -255 -229
rect -264 -231 -255 -230
rect -253 -231 -251 -229
rect -264 -234 -251 -231
rect -226 -229 -220 -225
rect -191 -223 -185 -222
rect -191 -225 -189 -223
rect -187 -225 -185 -223
rect -191 -229 -185 -225
rect -226 -230 -217 -229
rect -226 -232 -224 -230
rect -222 -232 -217 -230
rect -226 -233 -217 -232
rect -191 -230 -182 -229
rect -191 -232 -189 -230
rect -187 -232 -182 -230
rect -191 -233 -182 -232
rect -363 -252 -362 -250
rect -360 -252 -359 -250
rect -363 -256 -359 -252
rect -361 -258 -359 -256
rect -363 -267 -359 -258
rect -350 -247 -344 -246
rect -350 -249 -348 -247
rect -346 -249 -344 -247
rect -350 -253 -344 -249
rect -333 -247 -320 -246
rect -333 -249 -326 -247
rect -324 -249 -320 -247
rect -333 -250 -320 -249
rect -350 -256 -337 -253
rect -350 -258 -349 -256
rect -347 -258 -337 -256
rect -350 -259 -337 -258
rect -333 -254 -329 -250
rect -333 -256 -332 -254
rect -330 -256 -329 -254
rect -309 -249 -305 -238
rect -296 -239 -274 -238
rect -296 -241 -287 -239
rect -285 -240 -274 -239
rect -285 -241 -282 -240
rect -296 -242 -282 -241
rect -280 -242 -274 -240
rect -255 -236 -251 -234
rect -253 -238 -251 -236
rect -309 -251 -308 -249
rect -306 -251 -305 -249
rect -333 -259 -329 -256
rect -309 -257 -305 -251
rect -307 -259 -305 -257
rect -296 -247 -290 -246
rect -296 -249 -294 -247
rect -292 -249 -290 -247
rect -296 -253 -290 -249
rect -279 -247 -266 -246
rect -279 -249 -272 -247
rect -270 -249 -266 -247
rect -279 -250 -266 -249
rect -296 -256 -283 -253
rect -296 -258 -295 -256
rect -293 -258 -283 -256
rect -296 -259 -283 -258
rect -279 -254 -275 -250
rect -279 -256 -278 -254
rect -276 -256 -275 -254
rect -255 -249 -251 -238
rect -237 -241 -233 -237
rect -237 -242 -225 -241
rect -237 -244 -228 -242
rect -226 -244 -225 -242
rect -237 -245 -225 -244
rect -255 -251 -254 -249
rect -252 -251 -251 -249
rect -279 -259 -275 -256
rect -309 -267 -305 -259
rect -255 -257 -251 -251
rect -245 -249 -241 -245
rect -229 -247 -225 -245
rect -229 -249 -228 -247
rect -226 -249 -225 -247
rect -245 -250 -233 -249
rect -245 -252 -244 -250
rect -242 -252 -238 -250
rect -236 -252 -233 -250
rect -229 -251 -225 -249
rect -245 -253 -233 -252
rect -253 -259 -251 -257
rect -237 -259 -233 -253
rect -221 -255 -217 -233
rect -202 -241 -198 -237
rect -202 -242 -190 -241
rect -202 -244 -197 -242
rect -195 -244 -190 -242
rect -202 -245 -190 -244
rect -210 -249 -206 -245
rect -194 -247 -190 -245
rect -194 -249 -193 -247
rect -191 -249 -190 -247
rect -210 -250 -198 -249
rect -210 -252 -209 -250
rect -207 -252 -203 -250
rect -201 -252 -198 -250
rect -194 -251 -190 -249
rect -210 -253 -198 -252
rect -221 -257 -220 -255
rect -218 -257 -217 -255
rect -255 -267 -251 -259
rect -221 -261 -217 -257
rect -202 -259 -198 -253
rect -186 -257 -182 -233
rect -162 -238 -156 -230
rect -130 -229 -125 -221
rect -130 -230 -129 -229
rect -138 -231 -129 -230
rect -127 -231 -125 -229
rect -138 -234 -125 -231
rect -170 -239 -148 -238
rect -170 -241 -161 -239
rect -159 -240 -148 -239
rect -159 -241 -156 -240
rect -170 -242 -156 -241
rect -154 -242 -148 -240
rect -129 -236 -125 -234
rect -112 -231 -100 -229
rect -112 -233 -104 -231
rect -102 -233 -100 -231
rect -112 -235 -100 -233
rect -86 -231 -74 -229
rect -86 -233 -78 -231
rect -76 -233 -74 -231
rect -86 -235 -74 -233
rect -127 -238 -125 -236
rect -186 -259 -185 -257
rect -183 -259 -182 -257
rect -170 -247 -164 -246
rect -170 -249 -168 -247
rect -166 -249 -164 -247
rect -170 -253 -164 -249
rect -153 -247 -140 -246
rect -153 -249 -146 -247
rect -144 -249 -140 -247
rect -153 -250 -140 -249
rect -170 -256 -157 -253
rect -170 -258 -169 -256
rect -167 -258 -157 -256
rect -170 -259 -157 -258
rect -153 -255 -149 -250
rect -129 -253 -125 -238
rect -104 -238 -100 -235
rect -102 -240 -100 -238
rect -120 -247 -108 -245
rect -120 -249 -118 -247
rect -116 -249 -111 -247
rect -109 -249 -108 -247
rect -120 -251 -108 -249
rect -129 -255 -128 -253
rect -126 -255 -125 -253
rect -153 -257 -152 -255
rect -150 -257 -149 -255
rect -153 -259 -149 -257
rect -229 -263 -217 -261
rect -234 -264 -217 -263
rect -234 -266 -232 -264
rect -230 -266 -217 -264
rect -234 -267 -217 -266
rect -186 -261 -182 -259
rect -194 -263 -182 -261
rect -129 -257 -125 -255
rect -127 -259 -125 -257
rect -199 -264 -182 -263
rect -199 -266 -197 -264
rect -195 -266 -182 -264
rect -199 -267 -182 -266
rect -129 -267 -125 -259
rect -112 -259 -108 -251
rect -104 -250 -100 -240
rect -78 -238 -74 -235
rect -57 -238 -51 -230
rect -25 -229 -20 -221
rect -25 -230 -24 -229
rect -33 -231 -24 -230
rect -22 -231 -20 -229
rect -33 -234 -20 -231
rect -76 -240 -74 -238
rect -104 -252 -103 -250
rect -101 -252 -100 -250
rect -94 -247 -82 -245
rect -94 -249 -93 -247
rect -91 -249 -85 -247
rect -83 -249 -82 -247
rect -94 -251 -82 -249
rect -104 -256 -100 -252
rect -102 -258 -100 -256
rect -104 -267 -100 -258
rect -86 -259 -82 -251
rect -78 -250 -74 -240
rect -65 -239 -43 -238
rect -65 -241 -56 -239
rect -54 -240 -43 -239
rect -54 -241 -51 -240
rect -65 -242 -51 -241
rect -49 -242 -43 -240
rect -24 -236 -20 -234
rect -22 -238 -20 -236
rect -3 -238 3 -230
rect 29 -229 34 -221
rect 99 -217 106 -216
rect 59 -223 65 -222
rect 59 -225 61 -223
rect 63 -225 65 -223
rect 29 -230 30 -229
rect 21 -231 30 -230
rect 32 -231 34 -229
rect 21 -234 34 -231
rect 59 -229 65 -225
rect 94 -223 100 -222
rect 94 -225 96 -223
rect 98 -225 100 -223
rect 94 -229 100 -225
rect 59 -230 68 -229
rect 59 -232 61 -230
rect 63 -232 68 -230
rect 59 -233 68 -232
rect 94 -230 103 -229
rect 94 -232 96 -230
rect 98 -232 103 -230
rect 94 -233 103 -232
rect -78 -252 -77 -250
rect -75 -252 -74 -250
rect -78 -256 -74 -252
rect -76 -258 -74 -256
rect -78 -267 -74 -258
rect -65 -247 -59 -246
rect -65 -249 -63 -247
rect -61 -249 -59 -247
rect -65 -253 -59 -249
rect -48 -247 -35 -246
rect -48 -249 -41 -247
rect -39 -249 -35 -247
rect -48 -250 -35 -249
rect -65 -256 -52 -253
rect -65 -258 -64 -256
rect -62 -258 -52 -256
rect -65 -259 -52 -258
rect -48 -254 -44 -250
rect -48 -256 -47 -254
rect -45 -256 -44 -254
rect -24 -249 -20 -238
rect -11 -239 11 -238
rect -11 -241 -2 -239
rect 0 -240 11 -239
rect 0 -241 3 -240
rect -11 -242 3 -241
rect 5 -242 11 -240
rect 30 -236 34 -234
rect 32 -238 34 -236
rect -24 -251 -23 -249
rect -21 -251 -20 -249
rect -48 -259 -44 -256
rect -24 -257 -20 -251
rect -22 -259 -20 -257
rect -11 -247 -5 -246
rect -11 -249 -9 -247
rect -7 -249 -5 -247
rect -11 -253 -5 -249
rect 6 -247 19 -246
rect 6 -249 13 -247
rect 15 -249 19 -247
rect 6 -250 19 -249
rect -11 -256 2 -253
rect -11 -258 -10 -256
rect -8 -258 2 -256
rect -11 -259 2 -258
rect 6 -254 10 -250
rect 6 -256 7 -254
rect 9 -256 10 -254
rect 30 -249 34 -238
rect 48 -241 52 -237
rect 48 -242 60 -241
rect 48 -244 57 -242
rect 59 -244 60 -242
rect 48 -245 60 -244
rect 30 -251 31 -249
rect 33 -251 34 -249
rect 6 -259 10 -256
rect -24 -267 -20 -259
rect 30 -257 34 -251
rect 40 -249 44 -245
rect 56 -247 60 -245
rect 56 -249 57 -247
rect 59 -249 60 -247
rect 40 -250 52 -249
rect 40 -252 41 -250
rect 43 -252 47 -250
rect 49 -252 52 -250
rect 56 -251 60 -249
rect 40 -253 52 -252
rect 32 -259 34 -257
rect 48 -259 52 -253
rect 64 -255 68 -233
rect 83 -241 87 -237
rect 83 -242 95 -241
rect 83 -244 88 -242
rect 90 -244 95 -242
rect 83 -245 95 -244
rect 75 -249 79 -245
rect 91 -247 95 -245
rect 91 -249 92 -247
rect 94 -249 95 -247
rect 75 -250 87 -249
rect 75 -252 76 -250
rect 78 -252 82 -250
rect 84 -252 87 -250
rect 91 -251 95 -249
rect 75 -253 87 -252
rect 64 -257 65 -255
rect 67 -257 68 -255
rect 30 -267 34 -259
rect 64 -261 68 -257
rect 83 -259 87 -253
rect 99 -257 103 -233
rect 123 -238 129 -230
rect 155 -229 160 -221
rect 155 -230 156 -229
rect 147 -231 156 -230
rect 158 -231 160 -229
rect 147 -234 160 -231
rect 115 -239 137 -238
rect 115 -241 124 -239
rect 126 -240 137 -239
rect 126 -241 129 -240
rect 115 -242 129 -241
rect 131 -242 137 -240
rect 156 -236 160 -234
rect 173 -231 185 -229
rect 173 -233 181 -231
rect 183 -233 185 -231
rect 173 -235 185 -233
rect 199 -231 211 -229
rect 199 -233 207 -231
rect 209 -233 211 -231
rect 199 -235 211 -233
rect 158 -238 160 -236
rect 99 -259 100 -257
rect 102 -259 103 -257
rect 115 -247 121 -246
rect 115 -249 117 -247
rect 119 -249 121 -247
rect 115 -253 121 -249
rect 132 -247 145 -246
rect 132 -249 139 -247
rect 141 -249 145 -247
rect 132 -250 145 -249
rect 115 -256 128 -253
rect 115 -258 116 -256
rect 118 -258 128 -256
rect 115 -259 128 -258
rect 132 -255 136 -250
rect 156 -253 160 -238
rect 181 -238 185 -235
rect 183 -240 185 -238
rect 165 -247 177 -245
rect 165 -249 167 -247
rect 169 -249 174 -247
rect 176 -249 177 -247
rect 165 -251 177 -249
rect 156 -255 157 -253
rect 159 -255 160 -253
rect 132 -257 133 -255
rect 135 -257 136 -255
rect 132 -259 136 -257
rect 56 -263 68 -261
rect 51 -264 68 -263
rect 51 -266 53 -264
rect 55 -266 68 -264
rect 51 -267 68 -266
rect 99 -261 103 -259
rect 91 -263 103 -261
rect 156 -257 160 -255
rect 158 -259 160 -257
rect 86 -264 103 -263
rect 86 -266 88 -264
rect 90 -266 103 -264
rect 86 -267 103 -266
rect 156 -267 160 -259
rect 173 -259 177 -251
rect 181 -250 185 -240
rect 207 -238 211 -235
rect 228 -238 234 -230
rect 260 -229 265 -221
rect 260 -230 261 -229
rect 252 -231 261 -230
rect 263 -231 265 -229
rect 252 -234 265 -231
rect 209 -240 211 -238
rect 181 -252 182 -250
rect 184 -252 185 -250
rect 191 -247 203 -245
rect 191 -249 192 -247
rect 194 -249 200 -247
rect 202 -249 203 -247
rect 191 -251 203 -249
rect 181 -256 185 -252
rect 183 -258 185 -256
rect 181 -267 185 -258
rect 199 -259 203 -251
rect 207 -250 211 -240
rect 220 -239 242 -238
rect 220 -241 229 -239
rect 231 -240 242 -239
rect 231 -241 234 -240
rect 220 -242 234 -241
rect 236 -242 242 -240
rect 261 -236 265 -234
rect 263 -238 265 -236
rect 282 -238 288 -230
rect 314 -229 319 -221
rect 384 -217 391 -216
rect 344 -223 350 -222
rect 344 -225 346 -223
rect 348 -225 350 -223
rect 314 -230 315 -229
rect 306 -231 315 -230
rect 317 -231 319 -229
rect 306 -234 319 -231
rect 344 -229 350 -225
rect 379 -223 385 -222
rect 379 -225 381 -223
rect 383 -225 385 -223
rect 379 -229 385 -225
rect 344 -230 353 -229
rect 344 -232 346 -230
rect 348 -232 353 -230
rect 344 -233 353 -232
rect 379 -230 388 -229
rect 379 -232 381 -230
rect 383 -232 388 -230
rect 379 -233 388 -232
rect 207 -252 208 -250
rect 210 -252 211 -250
rect 207 -256 211 -252
rect 209 -258 211 -256
rect 207 -267 211 -258
rect 220 -247 226 -246
rect 220 -249 222 -247
rect 224 -249 226 -247
rect 220 -253 226 -249
rect 237 -247 250 -246
rect 237 -249 244 -247
rect 246 -249 250 -247
rect 237 -250 250 -249
rect 220 -256 233 -253
rect 220 -258 221 -256
rect 223 -258 233 -256
rect 220 -259 233 -258
rect 237 -254 241 -250
rect 237 -256 238 -254
rect 240 -256 241 -254
rect 261 -249 265 -238
rect 274 -239 296 -238
rect 274 -241 283 -239
rect 285 -240 296 -239
rect 285 -241 288 -240
rect 274 -242 288 -241
rect 290 -242 296 -240
rect 315 -236 319 -234
rect 317 -238 319 -236
rect 261 -251 262 -249
rect 264 -251 265 -249
rect 237 -259 241 -256
rect 261 -257 265 -251
rect 263 -259 265 -257
rect 274 -247 280 -246
rect 274 -249 276 -247
rect 278 -249 280 -247
rect 274 -253 280 -249
rect 291 -247 304 -246
rect 291 -249 298 -247
rect 300 -249 304 -247
rect 291 -250 304 -249
rect 274 -256 287 -253
rect 274 -258 275 -256
rect 277 -258 287 -256
rect 274 -259 287 -258
rect 291 -254 295 -250
rect 291 -256 292 -254
rect 294 -256 295 -254
rect 315 -249 319 -238
rect 333 -241 337 -237
rect 333 -242 345 -241
rect 333 -244 342 -242
rect 344 -244 345 -242
rect 333 -245 345 -244
rect 315 -251 316 -249
rect 318 -251 319 -249
rect 291 -259 295 -256
rect 261 -267 265 -259
rect 315 -257 319 -251
rect 325 -249 329 -245
rect 341 -247 345 -245
rect 341 -249 342 -247
rect 344 -249 345 -247
rect 325 -250 337 -249
rect 325 -252 326 -250
rect 328 -252 332 -250
rect 334 -252 337 -250
rect 341 -251 345 -249
rect 325 -253 337 -252
rect 317 -259 319 -257
rect 333 -259 337 -253
rect 349 -255 353 -233
rect 368 -241 372 -237
rect 368 -242 380 -241
rect 368 -244 373 -242
rect 375 -244 380 -242
rect 368 -245 380 -244
rect 360 -249 364 -245
rect 376 -247 380 -245
rect 376 -249 377 -247
rect 379 -249 380 -247
rect 360 -250 372 -249
rect 360 -252 361 -250
rect 363 -252 367 -250
rect 369 -252 372 -250
rect 376 -251 380 -249
rect 360 -253 372 -252
rect 349 -257 350 -255
rect 352 -257 353 -255
rect 315 -267 319 -259
rect 349 -261 353 -257
rect 368 -259 372 -253
rect 384 -257 388 -233
rect 408 -238 414 -230
rect 440 -229 445 -221
rect 440 -230 441 -229
rect 432 -231 441 -230
rect 443 -231 445 -229
rect 478 -230 482 -221
rect 432 -234 445 -231
rect 400 -239 422 -238
rect 400 -241 409 -239
rect 411 -240 422 -239
rect 411 -241 414 -240
rect 400 -242 414 -241
rect 416 -242 422 -240
rect 441 -236 445 -234
rect 443 -238 445 -236
rect 384 -259 385 -257
rect 387 -259 388 -257
rect 400 -247 406 -246
rect 400 -249 402 -247
rect 404 -249 406 -247
rect 400 -253 406 -249
rect 417 -247 430 -246
rect 417 -249 424 -247
rect 426 -249 430 -247
rect 417 -250 430 -249
rect 400 -256 413 -253
rect 400 -258 401 -256
rect 403 -258 413 -256
rect 400 -259 413 -258
rect 417 -255 421 -250
rect 441 -253 445 -238
rect 459 -234 522 -230
rect 459 -235 465 -234
rect 459 -237 460 -235
rect 462 -237 465 -235
rect 459 -239 465 -237
rect 459 -241 461 -239
rect 463 -241 465 -239
rect 459 -242 465 -241
rect 469 -240 475 -238
rect 469 -242 470 -240
rect 472 -242 475 -240
rect 485 -239 514 -238
rect 485 -241 487 -239
rect 489 -241 493 -239
rect 495 -241 514 -239
rect 485 -242 514 -241
rect 469 -245 475 -242
rect 469 -247 471 -245
rect 473 -246 475 -245
rect 473 -247 506 -246
rect 469 -250 506 -247
rect 441 -255 442 -253
rect 444 -255 445 -253
rect 502 -251 506 -250
rect 510 -251 514 -242
rect 518 -241 522 -234
rect 520 -243 522 -241
rect 518 -245 522 -243
rect 502 -253 503 -251
rect 505 -253 506 -251
rect 534 -231 538 -221
rect 570 -230 574 -221
rect 536 -233 538 -231
rect 534 -238 538 -233
rect 536 -240 538 -238
rect 417 -257 418 -255
rect 420 -257 421 -255
rect 417 -259 421 -257
rect 341 -263 353 -261
rect 336 -264 353 -263
rect 336 -266 338 -264
rect 340 -266 353 -264
rect 336 -267 353 -266
rect 384 -261 388 -259
rect 376 -263 388 -261
rect 441 -257 445 -255
rect 443 -259 445 -257
rect 475 -255 497 -254
rect 475 -257 477 -255
rect 479 -257 482 -255
rect 484 -257 493 -255
rect 495 -257 497 -255
rect 475 -258 497 -257
rect 371 -264 388 -263
rect 371 -266 373 -264
rect 375 -266 388 -264
rect 371 -267 388 -266
rect 441 -267 445 -259
rect 478 -267 482 -258
rect 502 -259 506 -253
rect 534 -262 538 -240
rect 551 -234 614 -230
rect 551 -235 557 -234
rect 551 -237 554 -235
rect 556 -237 557 -235
rect 551 -239 557 -237
rect 551 -241 553 -239
rect 555 -241 557 -239
rect 551 -242 557 -241
rect 561 -241 567 -238
rect 561 -243 562 -241
rect 564 -243 567 -241
rect 577 -239 606 -238
rect 577 -241 579 -239
rect 581 -241 599 -239
rect 601 -241 606 -239
rect 577 -242 606 -241
rect 561 -245 567 -243
rect 561 -247 563 -245
rect 565 -246 567 -245
rect 565 -247 598 -246
rect 561 -250 598 -247
rect 594 -251 598 -250
rect 602 -251 606 -242
rect 610 -241 614 -234
rect 612 -243 614 -241
rect 610 -245 614 -243
rect 594 -253 595 -251
rect 597 -253 598 -251
rect 626 -231 630 -221
rect 628 -233 630 -231
rect 626 -238 630 -233
rect 628 -240 630 -238
rect 567 -255 589 -254
rect 567 -257 569 -255
rect 571 -257 572 -255
rect 574 -257 585 -255
rect 587 -257 589 -255
rect 567 -258 589 -257
rect 524 -264 538 -262
rect 524 -266 534 -264
rect 536 -266 538 -264
rect 524 -267 538 -266
rect 570 -267 574 -258
rect 594 -259 598 -253
rect 626 -262 630 -240
rect 616 -264 630 -262
rect 616 -266 626 -264
rect 628 -266 630 -264
rect 616 -267 630 -266
rect -690 -273 744 -272
rect -690 -275 -687 -273
rect -685 -275 -675 -273
rect -673 -275 -661 -273
rect -659 -275 -649 -273
rect -647 -275 -605 -273
rect -603 -275 -595 -273
rect -593 -275 -551 -273
rect -549 -275 -541 -273
rect -539 -275 -527 -273
rect -525 -275 -506 -273
rect -504 -275 -492 -273
rect -490 -275 -471 -273
rect -469 -275 -425 -273
rect -423 -275 -415 -273
rect -413 -275 -402 -273
rect -400 -275 -390 -273
rect -388 -275 -376 -273
rect -374 -275 -364 -273
rect -362 -275 -320 -273
rect -318 -275 -310 -273
rect -308 -275 -266 -273
rect -264 -275 -256 -273
rect -254 -275 -242 -273
rect -240 -275 -221 -273
rect -219 -275 -207 -273
rect -205 -275 -186 -273
rect -184 -275 -140 -273
rect -138 -275 -130 -273
rect -128 -275 -117 -273
rect -115 -275 -105 -273
rect -103 -275 -91 -273
rect -89 -275 -79 -273
rect -77 -275 -35 -273
rect -33 -275 -25 -273
rect -23 -275 19 -273
rect 21 -275 29 -273
rect 31 -275 43 -273
rect 45 -275 64 -273
rect 66 -275 78 -273
rect 80 -275 99 -273
rect 101 -275 145 -273
rect 147 -275 155 -273
rect 157 -275 168 -273
rect 170 -275 180 -273
rect 182 -275 194 -273
rect 196 -275 206 -273
rect 208 -275 250 -273
rect 252 -275 260 -273
rect 262 -275 304 -273
rect 306 -275 314 -273
rect 316 -275 328 -273
rect 330 -275 349 -273
rect 351 -275 363 -273
rect 365 -275 384 -273
rect 386 -275 430 -273
rect 432 -275 440 -273
rect 442 -275 461 -273
rect 463 -275 469 -273
rect 471 -275 479 -273
rect 481 -275 501 -273
rect 503 -275 523 -273
rect 525 -275 553 -273
rect 555 -275 561 -273
rect 563 -275 571 -273
rect 573 -275 593 -273
rect 595 -275 615 -273
rect 617 -275 744 -273
rect -690 -277 739 -275
rect 741 -277 744 -275
rect -690 -280 744 -277
rect -674 -286 -631 -285
rect -674 -288 -673 -286
rect -671 -288 -634 -286
rect -632 -288 -631 -286
rect -674 -289 -631 -288
rect -540 -286 -526 -285
rect -540 -288 -539 -286
rect -537 -288 -529 -286
rect -527 -288 -526 -286
rect -540 -289 -526 -288
rect -506 -286 -491 -285
rect -506 -288 -505 -286
rect -503 -288 -494 -286
rect -492 -288 -491 -286
rect -506 -289 -491 -288
rect -483 -286 -479 -285
rect -483 -288 -482 -286
rect -480 -288 -479 -286
rect -483 -289 -479 -288
rect -389 -286 -346 -285
rect -389 -288 -388 -286
rect -386 -288 -349 -286
rect -347 -288 -346 -286
rect -389 -289 -346 -288
rect -255 -286 -241 -285
rect -255 -288 -254 -286
rect -252 -288 -244 -286
rect -242 -288 -241 -286
rect -255 -289 -241 -288
rect -221 -286 -206 -285
rect -221 -288 -220 -286
rect -218 -288 -209 -286
rect -207 -288 -206 -286
rect -221 -289 -206 -288
rect -198 -286 -194 -285
rect -198 -288 -197 -286
rect -195 -288 -194 -286
rect -198 -289 -194 -288
rect -104 -286 -61 -285
rect -104 -288 -103 -286
rect -101 -288 -64 -286
rect -62 -288 -61 -286
rect -104 -289 -61 -288
rect 30 -286 44 -285
rect 30 -288 31 -286
rect 33 -288 41 -286
rect 43 -288 44 -286
rect 30 -289 44 -288
rect 64 -286 79 -285
rect 64 -288 65 -286
rect 67 -288 76 -286
rect 78 -288 79 -286
rect 64 -289 79 -288
rect 87 -286 91 -285
rect 87 -288 88 -286
rect 90 -288 91 -286
rect 87 -289 91 -288
rect 181 -286 224 -285
rect 181 -288 182 -286
rect 184 -288 221 -286
rect 223 -288 224 -286
rect 181 -289 224 -288
rect 315 -286 329 -285
rect 315 -288 316 -286
rect 318 -288 326 -286
rect 328 -288 329 -286
rect 315 -289 329 -288
rect 349 -286 364 -285
rect 349 -288 350 -286
rect 352 -288 361 -286
rect 363 -288 364 -286
rect 349 -289 364 -288
rect 372 -286 376 -285
rect 372 -288 373 -286
rect 375 -288 376 -286
rect 372 -289 376 -288
rect 459 -287 684 -286
rect 459 -289 460 -287
rect 462 -289 681 -287
rect 683 -289 684 -287
rect 459 -290 684 -289
rect -689 -294 -577 -293
rect -689 -296 -688 -294
rect -686 -296 -580 -294
rect -578 -296 -577 -294
rect -689 -297 -577 -296
rect -514 -294 -451 -293
rect -514 -296 -513 -294
rect -511 -296 -470 -294
rect -468 -296 -454 -294
rect -452 -296 -451 -294
rect -514 -297 -451 -296
rect -404 -294 -292 -293
rect -404 -296 -403 -294
rect -401 -296 -295 -294
rect -293 -296 -292 -294
rect -404 -297 -292 -296
rect -229 -294 -166 -293
rect -229 -296 -228 -294
rect -226 -296 -185 -294
rect -183 -296 -169 -294
rect -167 -296 -166 -294
rect -229 -297 -166 -296
rect -119 -294 -7 -293
rect -119 -296 -118 -294
rect -116 -296 -10 -294
rect -8 -296 -7 -294
rect -119 -297 -7 -296
rect 56 -294 119 -293
rect 56 -296 57 -294
rect 59 -296 100 -294
rect 102 -296 116 -294
rect 118 -296 119 -294
rect 56 -297 119 -296
rect 166 -294 278 -293
rect 166 -296 167 -294
rect 169 -296 275 -294
rect 277 -296 278 -294
rect 166 -297 278 -296
rect 341 -294 404 -293
rect 341 -296 342 -294
rect 344 -296 385 -294
rect 387 -296 401 -294
rect 403 -296 404 -294
rect 341 -297 404 -296
rect 441 -295 557 -294
rect 441 -297 442 -295
rect 444 -297 554 -295
rect 556 -297 557 -295
rect 441 -298 557 -297
rect 561 -295 660 -294
rect 561 -297 562 -295
rect 564 -297 657 -295
rect 659 -297 660 -295
rect 561 -298 660 -297
rect -699 -302 -660 -301
rect -699 -304 -698 -302
rect -696 -304 -663 -302
rect -661 -304 -660 -302
rect -699 -305 -660 -304
rect -648 -302 -569 -301
rect -648 -304 -647 -302
rect -645 -304 -626 -302
rect -624 -304 -572 -302
rect -570 -304 -569 -302
rect -648 -305 -569 -304
rect -363 -302 -284 -301
rect -363 -304 -362 -302
rect -360 -304 -341 -302
rect -339 -304 -287 -302
rect -285 -304 -284 -302
rect -363 -305 -284 -304
rect -78 -302 1 -301
rect -78 -304 -77 -302
rect -75 -304 -56 -302
rect -54 -304 -2 -302
rect 0 -304 1 -302
rect -78 -305 1 -304
rect 207 -302 286 -301
rect 207 -304 208 -302
rect 210 -304 229 -302
rect 231 -304 283 -302
rect 285 -304 286 -302
rect 207 -305 286 -304
rect 469 -303 692 -302
rect 469 -305 470 -303
rect 472 -305 689 -303
rect 691 -305 692 -303
rect 469 -306 692 -305
rect -594 -310 -479 -309
rect -594 -312 -593 -310
rect -591 -312 -482 -310
rect -480 -312 -479 -310
rect -594 -313 -479 -312
rect -309 -310 -194 -309
rect -309 -312 -308 -310
rect -306 -312 -197 -310
rect -195 -312 -194 -310
rect -309 -313 -194 -312
rect -24 -310 91 -309
rect -24 -312 -23 -310
rect -21 -312 88 -310
rect 90 -312 91 -310
rect -24 -313 91 -312
rect 261 -310 376 -309
rect 261 -312 262 -310
rect 264 -312 373 -310
rect 375 -312 376 -310
rect 261 -313 376 -312
rect 481 -311 700 -310
rect 481 -313 482 -311
rect 484 -313 697 -311
rect 699 -313 700 -311
rect 481 -314 700 -313
rect -664 -318 -443 -317
rect -664 -320 -663 -318
rect -661 -320 -446 -318
rect -444 -320 -443 -318
rect -664 -321 -443 -320
rect -379 -318 -158 -317
rect -379 -320 -378 -318
rect -376 -320 -161 -318
rect -159 -320 -158 -318
rect -379 -321 -158 -320
rect -94 -318 127 -317
rect -94 -320 -93 -318
rect -91 -320 124 -318
rect 126 -320 127 -318
rect -94 -321 127 -320
rect 191 -318 412 -317
rect 191 -320 192 -318
rect 194 -320 409 -318
rect 411 -320 412 -318
rect 191 -321 412 -320
rect 571 -319 708 -318
rect 571 -321 572 -319
rect 574 -321 705 -319
rect 707 -321 708 -319
rect 571 -322 708 -321
rect -618 -326 -434 -325
rect -618 -328 -617 -326
rect -615 -328 -563 -326
rect -561 -328 -437 -326
rect -435 -328 -434 -326
rect -618 -329 -434 -328
rect -333 -326 -149 -325
rect -333 -328 -332 -326
rect -330 -328 -278 -326
rect -276 -328 -152 -326
rect -150 -328 -149 -326
rect -333 -329 -149 -328
rect -48 -326 136 -325
rect -48 -328 -47 -326
rect -45 -328 7 -326
rect 9 -328 133 -326
rect 135 -328 136 -326
rect -48 -329 136 -328
rect 156 -326 203 -325
rect 156 -328 157 -326
rect 159 -328 200 -326
rect 202 -328 203 -326
rect 156 -329 203 -328
rect 237 -326 421 -325
rect 237 -328 238 -326
rect 240 -328 292 -326
rect 294 -328 418 -326
rect 420 -328 421 -326
rect 237 -329 421 -328
rect 598 -327 716 -326
rect 598 -329 599 -327
rect 601 -329 713 -327
rect 715 -329 716 -327
rect 598 -330 716 -329
rect -618 -334 593 -333
rect -618 -336 -617 -334
rect -615 -336 -332 -334
rect -330 -336 -47 -334
rect -45 -336 238 -334
rect 240 -335 636 -334
rect 240 -336 633 -335
rect -618 -337 633 -336
rect 635 -337 636 -335
rect 589 -338 636 -337
rect -664 -342 195 -341
rect -664 -344 -663 -342
rect -661 -344 -378 -342
rect -376 -344 -93 -342
rect -91 -344 192 -342
rect 194 -344 195 -342
rect -664 -345 195 -344
rect 199 -342 496 -341
rect 199 -344 200 -342
rect 202 -344 493 -342
rect 495 -344 496 -342
rect 199 -345 496 -344
rect -707 -350 -400 -349
rect -707 -352 -706 -350
rect -704 -352 -403 -350
rect -401 -352 -400 -350
rect -707 -353 -400 -352
rect -129 -350 161 -349
rect -129 -352 -128 -350
rect -126 -352 158 -350
rect 160 -352 161 -350
rect -129 -353 161 -352
rect 166 -350 644 -349
rect 166 -352 167 -350
rect 169 -352 641 -350
rect 643 -352 644 -350
rect 166 -353 644 -352
rect -715 -358 -685 -357
rect -715 -360 -714 -358
rect -712 -360 -688 -358
rect -686 -360 -685 -358
rect -715 -361 -685 -360
rect -119 -358 652 -357
rect -119 -360 -118 -358
rect -116 -360 649 -358
rect 651 -360 652 -358
rect -119 -361 652 -360
rect -414 -367 668 -366
rect -414 -369 -413 -367
rect -411 -369 665 -367
rect 667 -369 668 -367
rect -414 -370 668 -369
rect 157 -375 676 -374
rect 157 -377 158 -375
rect 160 -377 673 -375
rect 675 -377 676 -375
rect 157 -378 676 -377
<< alu2 >>
rect 178 318 182 319
rect 178 316 179 318
rect 181 316 182 318
rect 149 310 153 311
rect 149 308 150 310
rect 152 308 153 310
rect -104 302 -100 303
rect -104 300 -103 302
rect -101 300 -100 302
rect -715 294 -711 295
rect -715 292 -714 294
rect -712 292 -711 294
rect -738 143 -724 150
rect -738 141 -733 143
rect -731 141 -724 143
rect -738 -207 -724 141
rect -738 -209 -733 -207
rect -731 -209 -724 -207
rect -738 -216 -724 -209
rect -715 -24 -711 292
rect -689 294 -685 295
rect -689 292 -688 294
rect -686 292 -685 294
rect -715 -26 -714 -24
rect -712 -26 -711 -24
rect -715 -40 -711 -26
rect -715 -42 -714 -40
rect -712 -42 -711 -40
rect -715 -358 -711 -42
rect -707 286 -703 287
rect -707 284 -706 286
rect -704 284 -703 286
rect -707 -8 -703 284
rect -707 -10 -706 -8
rect -704 -10 -703 -8
rect -707 -56 -703 -10
rect -707 -58 -706 -56
rect -704 -58 -703 -56
rect -707 -350 -703 -58
rect -699 238 -695 239
rect -699 236 -698 238
rect -696 236 -695 238
rect -699 48 -695 236
rect -689 230 -685 292
rect -414 294 -410 295
rect -414 292 -413 294
rect -411 292 -410 294
rect -689 228 -688 230
rect -686 228 -685 230
rect -689 183 -685 228
rect -664 278 -660 279
rect -664 276 -663 278
rect -661 276 -660 278
rect -664 254 -660 276
rect -664 252 -663 254
rect -661 252 -660 254
rect -664 238 -660 252
rect -618 270 -614 271
rect -618 268 -617 270
rect -615 268 -614 270
rect -618 262 -614 268
rect -618 260 -617 262
rect -615 260 -614 262
rect -664 236 -663 238
rect -661 236 -660 238
rect -674 222 -670 223
rect -674 220 -673 222
rect -671 220 -670 222
rect -674 186 -670 220
rect -674 184 -673 186
rect -671 184 -670 186
rect -674 183 -670 184
rect -664 183 -660 236
rect -648 238 -644 239
rect -648 236 -647 238
rect -645 236 -644 238
rect -648 186 -644 236
rect -627 238 -623 239
rect -627 236 -626 238
rect -624 236 -623 238
rect -635 222 -631 223
rect -635 220 -634 222
rect -632 220 -631 222
rect -635 192 -631 220
rect -635 190 -634 192
rect -632 190 -631 192
rect -635 189 -631 190
rect -648 184 -647 186
rect -645 184 -644 186
rect -648 183 -644 184
rect -689 181 -688 183
rect -686 181 -685 183
rect -689 180 -685 181
rect -664 181 -663 183
rect -661 181 -660 183
rect -664 179 -660 181
rect -627 175 -623 236
rect -618 190 -614 260
rect -564 262 -560 263
rect -564 260 -563 262
rect -561 260 -560 262
rect -618 188 -617 190
rect -615 188 -614 190
rect -618 187 -614 188
rect -594 246 -590 247
rect -594 244 -593 246
rect -591 244 -590 246
rect -594 185 -590 244
rect -573 238 -569 239
rect -573 236 -572 238
rect -570 236 -569 238
rect -581 230 -577 231
rect -581 228 -580 230
rect -578 228 -577 230
rect -581 192 -577 228
rect -581 190 -580 192
rect -578 190 -577 192
rect -581 189 -577 190
rect -594 183 -593 185
rect -591 183 -590 185
rect -594 182 -590 183
rect -627 173 -626 175
rect -624 173 -623 175
rect -627 172 -623 173
rect -573 175 -569 236
rect -564 190 -560 260
rect -438 262 -434 263
rect -438 260 -437 262
rect -435 260 -434 262
rect -447 254 -443 255
rect -447 252 -446 254
rect -444 252 -443 254
rect -483 246 -479 247
rect -483 244 -482 246
rect -480 244 -479 246
rect -514 230 -510 231
rect -514 228 -513 230
rect -511 228 -510 230
rect -564 188 -563 190
rect -561 188 -560 190
rect -564 187 -560 188
rect -540 222 -536 223
rect -540 220 -539 222
rect -537 220 -536 222
rect -540 185 -536 220
rect -540 183 -539 185
rect -537 183 -536 185
rect -530 222 -526 223
rect -530 220 -529 222
rect -527 220 -526 222
rect -530 186 -526 220
rect -530 184 -529 186
rect -527 184 -526 186
rect -530 183 -526 184
rect -540 182 -536 183
rect -514 178 -510 228
rect -506 222 -502 223
rect -506 220 -505 222
rect -503 220 -502 222
rect -506 191 -502 220
rect -506 189 -505 191
rect -503 189 -502 191
rect -506 188 -502 189
rect -495 222 -491 223
rect -495 220 -494 222
rect -492 220 -491 222
rect -495 186 -491 220
rect -495 184 -494 186
rect -492 184 -491 186
rect -495 183 -491 184
rect -483 222 -479 244
rect -483 220 -482 222
rect -480 220 -479 222
rect -514 176 -513 178
rect -511 176 -510 178
rect -514 175 -510 176
rect -483 178 -479 220
rect -471 230 -467 231
rect -471 228 -470 230
rect -468 228 -467 230
rect -471 193 -467 228
rect -471 191 -470 193
rect -468 191 -467 193
rect -471 190 -467 191
rect -455 230 -451 231
rect -455 228 -454 230
rect -452 228 -451 230
rect -455 192 -451 228
rect -455 190 -454 192
rect -452 190 -451 192
rect -455 189 -451 190
rect -483 176 -482 178
rect -480 176 -479 178
rect -483 175 -479 176
rect -447 175 -443 252
rect -438 191 -434 260
rect -438 189 -437 191
rect -435 189 -434 191
rect -438 187 -434 189
rect -428 180 -424 214
rect -414 189 -410 292
rect -127 294 -123 295
rect -127 292 -126 294
rect -124 292 -123 294
rect -414 187 -413 189
rect -411 187 -410 189
rect -414 186 -410 187
rect -404 286 -400 287
rect -404 284 -403 286
rect -401 284 -400 286
rect -404 230 -400 284
rect -127 286 -123 292
rect -127 284 -126 286
rect -124 284 -123 286
rect -127 283 -123 284
rect -119 294 -115 295
rect -119 292 -118 294
rect -116 292 -115 294
rect -404 228 -403 230
rect -401 228 -400 230
rect -404 183 -400 228
rect -379 278 -375 279
rect -379 276 -378 278
rect -376 276 -375 278
rect -379 254 -375 276
rect -379 252 -378 254
rect -376 252 -375 254
rect -389 222 -385 223
rect -389 220 -388 222
rect -386 220 -385 222
rect -389 186 -385 220
rect -389 184 -388 186
rect -386 184 -385 186
rect -389 183 -385 184
rect -379 183 -375 252
rect -333 270 -329 271
rect -333 268 -332 270
rect -330 268 -329 270
rect -333 262 -329 268
rect -333 260 -332 262
rect -330 260 -329 262
rect -363 238 -359 239
rect -363 236 -362 238
rect -360 236 -359 238
rect -363 186 -359 236
rect -342 238 -338 239
rect -342 236 -341 238
rect -339 236 -338 238
rect -350 222 -346 223
rect -350 220 -349 222
rect -347 220 -346 222
rect -350 192 -346 220
rect -350 190 -349 192
rect -347 190 -346 192
rect -350 189 -346 190
rect -363 184 -362 186
rect -360 184 -359 186
rect -363 183 -359 184
rect -404 181 -403 183
rect -401 181 -400 183
rect -404 180 -400 181
rect -379 181 -378 183
rect -376 181 -375 183
rect -379 179 -375 181
rect -573 173 -572 175
rect -570 173 -569 175
rect -573 172 -569 173
rect -447 173 -446 175
rect -444 173 -443 175
rect -447 172 -443 173
rect -342 175 -338 236
rect -333 190 -329 260
rect -279 262 -275 263
rect -279 260 -278 262
rect -276 260 -275 262
rect -333 188 -332 190
rect -330 188 -329 190
rect -333 187 -329 188
rect -309 246 -305 247
rect -309 244 -308 246
rect -306 244 -305 246
rect -309 185 -305 244
rect -288 238 -284 239
rect -288 236 -287 238
rect -285 236 -284 238
rect -296 230 -292 231
rect -296 228 -295 230
rect -293 228 -292 230
rect -296 192 -292 228
rect -296 190 -295 192
rect -293 190 -292 192
rect -296 189 -292 190
rect -309 183 -308 185
rect -306 183 -305 185
rect -309 182 -305 183
rect -342 173 -341 175
rect -339 173 -338 175
rect -342 172 -338 173
rect -288 175 -284 236
rect -279 190 -275 260
rect -153 262 -149 263
rect -153 260 -152 262
rect -150 260 -149 262
rect -162 254 -158 255
rect -162 252 -161 254
rect -159 252 -158 254
rect -198 246 -194 247
rect -198 244 -197 246
rect -195 244 -194 246
rect -229 230 -225 231
rect -229 228 -228 230
rect -226 228 -225 230
rect -279 188 -278 190
rect -276 188 -275 190
rect -279 187 -275 188
rect -255 222 -251 223
rect -255 220 -254 222
rect -252 220 -251 222
rect -255 185 -251 220
rect -255 183 -254 185
rect -252 183 -251 185
rect -245 222 -241 223
rect -245 220 -244 222
rect -242 220 -241 222
rect -245 186 -241 220
rect -245 184 -244 186
rect -242 184 -241 186
rect -245 183 -241 184
rect -255 182 -251 183
rect -229 178 -225 228
rect -221 222 -217 223
rect -221 220 -220 222
rect -218 220 -217 222
rect -221 191 -217 220
rect -221 189 -220 191
rect -218 189 -217 191
rect -221 188 -217 189
rect -210 222 -206 223
rect -210 220 -209 222
rect -207 220 -206 222
rect -210 186 -206 220
rect -210 184 -209 186
rect -207 184 -206 186
rect -210 183 -206 184
rect -198 222 -194 244
rect -198 220 -197 222
rect -195 220 -194 222
rect -229 176 -228 178
rect -226 176 -225 178
rect -229 175 -225 176
rect -198 178 -194 220
rect -186 230 -182 231
rect -186 228 -185 230
rect -183 228 -182 230
rect -186 193 -182 228
rect -186 191 -185 193
rect -183 191 -182 193
rect -186 190 -182 191
rect -170 230 -166 231
rect -170 228 -169 230
rect -167 228 -166 230
rect -170 192 -166 228
rect -170 190 -169 192
rect -167 190 -166 192
rect -170 189 -166 190
rect -198 176 -197 178
rect -195 176 -194 178
rect -198 175 -194 176
rect -162 175 -158 252
rect -153 191 -149 260
rect -129 238 -125 239
rect -129 236 -128 238
rect -126 236 -125 238
rect -153 189 -152 191
rect -150 189 -149 191
rect -153 187 -149 189
rect -143 180 -139 214
rect -129 189 -125 236
rect -129 187 -128 189
rect -126 187 -125 189
rect -129 186 -125 187
rect -119 230 -115 292
rect -104 238 -100 300
rect 149 302 153 308
rect 149 300 150 302
rect 152 300 153 302
rect 149 299 153 300
rect 157 302 161 303
rect 157 300 158 302
rect 160 300 161 302
rect 157 286 161 300
rect 157 284 158 286
rect 160 284 161 286
rect 157 283 161 284
rect 166 286 170 287
rect 166 284 167 286
rect 169 284 170 286
rect -104 236 -103 238
rect -101 236 -100 238
rect -104 235 -100 236
rect -94 278 -90 279
rect -94 276 -93 278
rect -91 276 -90 278
rect -94 254 -90 276
rect -94 252 -93 254
rect -91 252 -90 254
rect -119 228 -118 230
rect -116 228 -115 230
rect -119 183 -115 228
rect -104 222 -100 223
rect -104 220 -103 222
rect -101 220 -100 222
rect -104 186 -100 220
rect -104 184 -103 186
rect -101 184 -100 186
rect -104 183 -100 184
rect -94 183 -90 252
rect -48 270 -44 271
rect -48 268 -47 270
rect -45 268 -44 270
rect -48 262 -44 268
rect -48 260 -47 262
rect -45 260 -44 262
rect -78 238 -74 239
rect -78 236 -77 238
rect -75 236 -74 238
rect -78 186 -74 236
rect -57 238 -53 239
rect -57 236 -56 238
rect -54 236 -53 238
rect -65 222 -61 223
rect -65 220 -64 222
rect -62 220 -61 222
rect -65 192 -61 220
rect -65 190 -64 192
rect -62 190 -61 192
rect -65 189 -61 190
rect -78 184 -77 186
rect -75 184 -74 186
rect -78 183 -74 184
rect -119 181 -118 183
rect -116 181 -115 183
rect -119 180 -115 181
rect -94 181 -93 183
rect -91 181 -90 183
rect -94 179 -90 181
rect -288 173 -287 175
rect -285 173 -284 175
rect -288 172 -284 173
rect -162 173 -161 175
rect -159 173 -158 175
rect -162 172 -158 173
rect -57 175 -53 236
rect -48 190 -44 260
rect 6 262 10 263
rect 6 260 7 262
rect 9 260 10 262
rect -48 188 -47 190
rect -45 188 -44 190
rect -48 187 -44 188
rect -24 246 -20 247
rect -24 244 -23 246
rect -21 244 -20 246
rect -24 185 -20 244
rect -3 238 1 239
rect -3 236 -2 238
rect 0 236 1 238
rect -11 230 -7 231
rect -11 228 -10 230
rect -8 228 -7 230
rect -11 192 -7 228
rect -11 190 -10 192
rect -8 190 -7 192
rect -11 189 -7 190
rect -24 183 -23 185
rect -21 183 -20 185
rect -24 182 -20 183
rect -57 173 -56 175
rect -54 173 -53 175
rect -57 172 -53 173
rect -3 175 1 236
rect 6 190 10 260
rect 132 262 136 263
rect 132 260 133 262
rect 135 260 136 262
rect 123 254 127 255
rect 123 252 124 254
rect 126 252 127 254
rect 87 246 91 247
rect 87 244 88 246
rect 90 244 91 246
rect 56 230 60 231
rect 56 228 57 230
rect 59 228 60 230
rect 6 188 7 190
rect 9 188 10 190
rect 6 187 10 188
rect 30 222 34 223
rect 30 220 31 222
rect 33 220 34 222
rect 30 185 34 220
rect 30 183 31 185
rect 33 183 34 185
rect 40 222 44 223
rect 40 220 41 222
rect 43 220 44 222
rect 40 186 44 220
rect 40 184 41 186
rect 43 184 44 186
rect 40 183 44 184
rect 30 182 34 183
rect 56 178 60 228
rect 64 222 68 223
rect 64 220 65 222
rect 67 220 68 222
rect 64 191 68 220
rect 64 189 65 191
rect 67 189 68 191
rect 64 188 68 189
rect 75 222 79 223
rect 75 220 76 222
rect 78 220 79 222
rect 75 186 79 220
rect 75 184 76 186
rect 78 184 79 186
rect 75 183 79 184
rect 87 222 91 244
rect 87 220 88 222
rect 90 220 91 222
rect 56 176 57 178
rect 59 176 60 178
rect 56 175 60 176
rect 87 178 91 220
rect 99 230 103 231
rect 99 228 100 230
rect 102 228 103 230
rect 99 193 103 228
rect 99 191 100 193
rect 102 191 103 193
rect 99 190 103 191
rect 115 230 119 231
rect 115 228 116 230
rect 118 228 119 230
rect 115 192 119 228
rect 115 190 116 192
rect 118 190 119 192
rect 115 189 119 190
rect 87 176 88 178
rect 90 176 91 178
rect 87 175 91 176
rect 123 175 127 252
rect 132 191 136 260
rect 156 242 160 243
rect 156 240 157 242
rect 159 240 160 242
rect 132 189 133 191
rect 135 189 136 191
rect 132 187 136 189
rect 142 180 146 214
rect 156 189 160 240
rect 156 187 157 189
rect 159 187 160 189
rect 156 186 160 187
rect 166 230 170 284
rect 178 242 182 316
rect 672 318 676 319
rect 672 316 673 318
rect 675 316 676 318
rect 664 310 668 311
rect 664 308 665 310
rect 667 308 668 310
rect 656 302 660 303
rect 656 300 657 302
rect 659 300 660 302
rect 648 294 652 295
rect 648 292 649 294
rect 651 292 652 294
rect 640 286 644 287
rect 640 284 641 286
rect 643 284 644 286
rect 178 240 179 242
rect 181 240 182 242
rect 178 239 182 240
rect 191 278 195 279
rect 191 276 192 278
rect 194 276 195 278
rect 191 254 195 276
rect 441 278 445 279
rect 441 276 442 278
rect 444 276 445 278
rect 191 252 192 254
rect 194 252 195 254
rect 166 228 167 230
rect 169 228 170 230
rect 166 183 170 228
rect 181 222 185 223
rect 181 220 182 222
rect 184 220 185 222
rect 181 186 185 220
rect 181 184 182 186
rect 184 184 185 186
rect 181 183 185 184
rect 191 183 195 252
rect 237 270 241 271
rect 237 268 238 270
rect 240 268 241 270
rect 237 262 241 268
rect 237 260 238 262
rect 240 260 241 262
rect 207 238 211 239
rect 207 236 208 238
rect 210 236 211 238
rect 207 186 211 236
rect 228 238 232 239
rect 228 236 229 238
rect 231 236 232 238
rect 220 222 224 223
rect 220 220 221 222
rect 223 220 224 222
rect 220 192 224 220
rect 220 190 221 192
rect 223 190 224 192
rect 220 189 224 190
rect 207 184 208 186
rect 210 184 211 186
rect 207 183 211 184
rect 166 181 167 183
rect 169 181 170 183
rect 166 180 170 181
rect 191 181 192 183
rect 194 181 195 183
rect 191 179 195 181
rect -3 173 -2 175
rect 0 173 1 175
rect -3 172 1 173
rect 123 173 124 175
rect 126 173 127 175
rect 123 172 127 173
rect 228 175 232 236
rect 237 190 241 260
rect 291 262 295 263
rect 291 260 292 262
rect 294 260 295 262
rect 237 188 238 190
rect 240 188 241 190
rect 237 187 241 188
rect 261 246 265 247
rect 261 244 262 246
rect 264 244 265 246
rect 261 185 265 244
rect 282 238 286 239
rect 282 236 283 238
rect 285 236 286 238
rect 274 230 278 231
rect 274 228 275 230
rect 277 228 278 230
rect 274 192 278 228
rect 274 190 275 192
rect 277 190 278 192
rect 274 189 278 190
rect 261 183 262 185
rect 264 183 265 185
rect 261 182 265 183
rect 228 173 229 175
rect 231 173 232 175
rect 228 172 232 173
rect 282 175 286 236
rect 291 190 295 260
rect 417 262 421 263
rect 417 260 418 262
rect 420 260 421 262
rect 408 254 412 255
rect 408 252 409 254
rect 411 252 412 254
rect 372 246 376 247
rect 372 244 373 246
rect 375 244 376 246
rect 341 230 345 231
rect 341 228 342 230
rect 344 228 345 230
rect 291 188 292 190
rect 294 188 295 190
rect 291 187 295 188
rect 315 222 319 223
rect 315 220 316 222
rect 318 220 319 222
rect 315 185 319 220
rect 315 183 316 185
rect 318 183 319 185
rect 325 222 329 223
rect 325 220 326 222
rect 328 220 329 222
rect 325 186 329 220
rect 325 184 326 186
rect 328 184 329 186
rect 325 183 329 184
rect 315 182 319 183
rect 341 178 345 228
rect 349 222 353 223
rect 349 220 350 222
rect 352 220 353 222
rect 349 191 353 220
rect 349 189 350 191
rect 352 189 353 191
rect 349 188 353 189
rect 360 222 364 223
rect 360 220 361 222
rect 363 220 364 222
rect 360 186 364 220
rect 360 184 361 186
rect 363 184 364 186
rect 360 183 364 184
rect 372 222 376 244
rect 372 220 373 222
rect 375 220 376 222
rect 341 176 342 178
rect 344 176 345 178
rect 341 175 345 176
rect 372 178 376 220
rect 384 230 388 231
rect 384 228 385 230
rect 387 228 388 230
rect 384 193 388 228
rect 384 191 385 193
rect 387 191 388 193
rect 384 190 388 191
rect 400 230 404 231
rect 400 228 401 230
rect 403 228 404 230
rect 400 192 404 228
rect 400 190 401 192
rect 403 190 404 192
rect 400 189 404 190
rect 372 176 373 178
rect 375 176 376 178
rect 372 175 376 176
rect 408 175 412 252
rect 417 191 421 260
rect 417 189 418 191
rect 420 189 421 191
rect 417 187 421 189
rect 427 180 431 214
rect 441 189 445 276
rect 514 270 518 271
rect 514 268 515 270
rect 517 268 518 270
rect 441 187 442 189
rect 444 187 445 189
rect 441 186 445 187
rect 454 262 458 263
rect 454 260 455 262
rect 457 260 458 262
rect 454 254 458 260
rect 454 252 455 254
rect 457 252 458 254
rect 454 187 458 252
rect 514 254 518 268
rect 514 252 515 254
rect 517 252 518 254
rect 478 246 482 247
rect 478 244 479 246
rect 481 244 482 246
rect 478 192 482 244
rect 478 190 479 192
rect 481 190 482 192
rect 478 189 482 190
rect 488 230 492 231
rect 488 228 489 230
rect 491 228 492 230
rect 454 185 455 187
rect 457 185 458 187
rect 454 184 458 185
rect 282 173 283 175
rect 285 173 286 175
rect 282 172 286 173
rect 408 173 409 175
rect 411 173 412 175
rect 408 172 412 173
rect 488 175 492 228
rect 499 222 503 223
rect 499 220 500 222
rect 502 220 503 222
rect 499 206 503 220
rect 499 191 504 206
rect 496 190 504 191
rect 496 188 497 190
rect 499 188 504 190
rect 496 187 504 188
rect 514 187 518 252
rect 632 262 636 263
rect 632 260 633 262
rect 635 260 636 262
rect 538 246 542 247
rect 538 244 539 246
rect 541 244 542 246
rect 538 192 542 244
rect 608 246 612 247
rect 608 244 609 246
rect 611 244 612 246
rect 538 190 539 192
rect 541 190 542 192
rect 538 189 542 190
rect 550 238 554 239
rect 550 236 551 238
rect 553 236 554 238
rect 550 192 554 236
rect 580 238 584 239
rect 580 236 581 238
rect 583 236 584 238
rect 550 190 551 192
rect 553 190 554 192
rect 550 189 554 190
rect 559 222 563 223
rect 559 220 560 222
rect 562 220 563 222
rect 559 189 563 220
rect 580 199 584 236
rect 580 197 581 199
rect 583 197 584 199
rect 580 195 584 197
rect 596 230 600 231
rect 596 228 597 230
rect 599 228 600 230
rect 514 185 515 187
rect 517 185 518 187
rect 514 184 518 185
rect 488 173 489 175
rect 491 173 492 175
rect 488 172 492 173
rect 559 175 568 189
rect 596 183 600 228
rect 596 181 597 183
rect 599 181 600 183
rect 596 179 600 181
rect 559 173 560 175
rect 562 173 568 175
rect 559 172 568 173
rect -627 111 -623 112
rect -627 109 -626 111
rect -624 109 -623 111
rect -699 46 -698 48
rect -696 46 -695 48
rect -699 -112 -695 46
rect -689 103 -685 104
rect -689 101 -688 103
rect -686 101 -685 103
rect -664 103 -660 105
rect -664 101 -663 103
rect -661 101 -660 103
rect -689 56 -685 101
rect -674 100 -670 101
rect -674 98 -673 100
rect -671 98 -670 100
rect -674 64 -670 98
rect -674 62 -673 64
rect -671 62 -670 64
rect -674 61 -670 62
rect -689 54 -688 56
rect -686 54 -685 56
rect -689 -24 -685 54
rect -664 48 -660 101
rect -664 46 -663 48
rect -661 46 -660 48
rect -664 32 -660 46
rect -648 100 -644 101
rect -648 98 -647 100
rect -645 98 -644 100
rect -648 48 -644 98
rect -635 94 -631 95
rect -635 92 -634 94
rect -632 92 -631 94
rect -635 64 -631 92
rect -635 62 -634 64
rect -632 62 -631 64
rect -635 61 -631 62
rect -648 46 -647 48
rect -645 46 -644 48
rect -648 45 -644 46
rect -627 48 -623 109
rect -573 111 -569 112
rect -573 109 -572 111
rect -570 109 -569 111
rect -447 111 -443 112
rect -447 109 -446 111
rect -444 109 -443 111
rect -594 101 -590 102
rect -594 99 -593 101
rect -591 99 -590 101
rect -627 46 -626 48
rect -624 46 -623 48
rect -627 45 -623 46
rect -618 96 -614 97
rect -618 94 -617 96
rect -615 94 -614 96
rect -664 30 -663 32
rect -661 30 -660 32
rect -664 8 -660 30
rect -618 24 -614 94
rect -594 40 -590 99
rect -581 94 -577 95
rect -581 92 -580 94
rect -578 92 -577 94
rect -581 56 -577 92
rect -581 54 -580 56
rect -578 54 -577 56
rect -581 53 -577 54
rect -573 48 -569 109
rect -514 108 -510 109
rect -514 106 -513 108
rect -511 106 -510 108
rect -540 101 -536 102
rect -540 99 -539 101
rect -537 99 -536 101
rect -573 46 -572 48
rect -570 46 -569 48
rect -573 45 -569 46
rect -564 96 -560 97
rect -564 94 -563 96
rect -561 94 -560 96
rect -594 38 -593 40
rect -591 38 -590 40
rect -594 37 -590 38
rect -618 22 -617 24
rect -615 22 -614 24
rect -618 16 -614 22
rect -564 24 -560 94
rect -540 64 -536 99
rect -540 62 -539 64
rect -537 62 -536 64
rect -540 61 -536 62
rect -530 100 -526 101
rect -530 98 -529 100
rect -527 98 -526 100
rect -530 64 -526 98
rect -530 62 -529 64
rect -527 62 -526 64
rect -530 61 -526 62
rect -514 56 -510 106
rect -483 108 -479 109
rect -483 106 -482 108
rect -480 106 -479 108
rect -495 100 -491 101
rect -495 98 -494 100
rect -492 98 -491 100
rect -506 95 -502 96
rect -506 93 -505 95
rect -503 93 -502 95
rect -506 64 -502 93
rect -506 62 -505 64
rect -503 62 -502 64
rect -506 61 -502 62
rect -495 64 -491 98
rect -495 62 -494 64
rect -492 62 -491 64
rect -495 61 -491 62
rect -483 64 -479 106
rect -455 94 -451 95
rect -483 62 -482 64
rect -480 62 -479 64
rect -514 54 -513 56
rect -511 54 -510 56
rect -514 53 -510 54
rect -483 40 -479 62
rect -471 93 -467 94
rect -471 91 -470 93
rect -468 91 -467 93
rect -471 56 -467 91
rect -471 54 -470 56
rect -468 54 -467 56
rect -471 53 -467 54
rect -455 92 -454 94
rect -452 92 -451 94
rect -455 56 -451 92
rect -455 54 -454 56
rect -452 54 -451 56
rect -455 53 -451 54
rect -483 38 -482 40
rect -480 38 -479 40
rect -483 37 -479 38
rect -447 32 -443 109
rect -342 111 -338 112
rect -342 109 -341 111
rect -339 109 -338 111
rect -447 30 -446 32
rect -444 30 -443 32
rect -447 29 -443 30
rect -438 95 -434 97
rect -438 93 -437 95
rect -435 93 -434 95
rect -564 22 -563 24
rect -561 22 -560 24
rect -564 21 -560 22
rect -438 24 -434 93
rect -428 70 -424 104
rect -404 103 -400 104
rect -404 101 -403 103
rect -401 101 -400 103
rect -379 103 -375 105
rect -379 101 -378 103
rect -376 101 -375 103
rect -414 97 -410 98
rect -414 95 -413 97
rect -411 95 -410 97
rect -438 22 -437 24
rect -435 22 -434 24
rect -438 21 -434 22
rect -618 14 -617 16
rect -615 14 -614 16
rect -618 13 -614 14
rect -664 6 -663 8
rect -661 6 -660 8
rect -664 5 -660 6
rect -414 0 -410 95
rect -414 -2 -413 0
rect -411 -2 -410 0
rect -414 -3 -410 -2
rect -404 56 -400 101
rect -389 100 -385 101
rect -389 98 -388 100
rect -386 98 -385 100
rect -389 64 -385 98
rect -389 62 -388 64
rect -386 62 -385 64
rect -389 61 -385 62
rect -404 54 -403 56
rect -401 54 -400 56
rect -404 -8 -400 54
rect -379 32 -375 101
rect -363 100 -359 101
rect -363 98 -362 100
rect -360 98 -359 100
rect -363 48 -359 98
rect -350 94 -346 95
rect -350 92 -349 94
rect -347 92 -346 94
rect -350 64 -346 92
rect -350 62 -349 64
rect -347 62 -346 64
rect -350 61 -346 62
rect -363 46 -362 48
rect -360 46 -359 48
rect -363 45 -359 46
rect -342 48 -338 109
rect -288 111 -284 112
rect -288 109 -287 111
rect -285 109 -284 111
rect -162 111 -158 112
rect -162 109 -161 111
rect -159 109 -158 111
rect -309 101 -305 102
rect -309 99 -308 101
rect -306 99 -305 101
rect -342 46 -341 48
rect -339 46 -338 48
rect -342 45 -338 46
rect -333 96 -329 97
rect -333 94 -332 96
rect -330 94 -329 96
rect -379 30 -378 32
rect -376 30 -375 32
rect -379 8 -375 30
rect -333 24 -329 94
rect -309 40 -305 99
rect -296 94 -292 95
rect -296 92 -295 94
rect -293 92 -292 94
rect -296 56 -292 92
rect -296 54 -295 56
rect -293 54 -292 56
rect -296 53 -292 54
rect -288 48 -284 109
rect -229 108 -225 109
rect -229 106 -228 108
rect -226 106 -225 108
rect -255 101 -251 102
rect -255 99 -254 101
rect -252 99 -251 101
rect -288 46 -287 48
rect -285 46 -284 48
rect -288 45 -284 46
rect -279 96 -275 97
rect -279 94 -278 96
rect -276 94 -275 96
rect -309 38 -308 40
rect -306 38 -305 40
rect -309 37 -305 38
rect -333 22 -332 24
rect -330 22 -329 24
rect -333 16 -329 22
rect -279 24 -275 94
rect -255 64 -251 99
rect -255 62 -254 64
rect -252 62 -251 64
rect -255 61 -251 62
rect -245 100 -241 101
rect -245 98 -244 100
rect -242 98 -241 100
rect -245 64 -241 98
rect -245 62 -244 64
rect -242 62 -241 64
rect -245 61 -241 62
rect -229 56 -225 106
rect -198 108 -194 109
rect -198 106 -197 108
rect -195 106 -194 108
rect -210 100 -206 101
rect -210 98 -209 100
rect -207 98 -206 100
rect -221 95 -217 96
rect -221 93 -220 95
rect -218 93 -217 95
rect -221 64 -217 93
rect -221 62 -220 64
rect -218 62 -217 64
rect -221 61 -217 62
rect -210 64 -206 98
rect -210 62 -209 64
rect -207 62 -206 64
rect -210 61 -206 62
rect -198 64 -194 106
rect -170 94 -166 95
rect -198 62 -197 64
rect -195 62 -194 64
rect -229 54 -228 56
rect -226 54 -225 56
rect -229 53 -225 54
rect -198 40 -194 62
rect -186 93 -182 94
rect -186 91 -185 93
rect -183 91 -182 93
rect -186 56 -182 91
rect -186 54 -185 56
rect -183 54 -182 56
rect -186 53 -182 54
rect -170 92 -169 94
rect -167 92 -166 94
rect -170 56 -166 92
rect -170 54 -169 56
rect -167 54 -166 56
rect -170 53 -166 54
rect -198 38 -197 40
rect -195 38 -194 40
rect -198 37 -194 38
rect -162 32 -158 109
rect -57 111 -53 112
rect -57 109 -56 111
rect -54 109 -53 111
rect -162 30 -161 32
rect -159 30 -158 32
rect -162 29 -158 30
rect -153 95 -149 97
rect -153 93 -152 95
rect -150 93 -149 95
rect -279 22 -278 24
rect -276 22 -275 24
rect -279 21 -275 22
rect -153 24 -149 93
rect -143 70 -139 104
rect -119 103 -115 104
rect -119 101 -118 103
rect -116 101 -115 103
rect -94 103 -90 105
rect -94 101 -93 103
rect -91 101 -90 103
rect -129 97 -125 98
rect -129 95 -128 97
rect -126 95 -125 97
rect -153 22 -152 24
rect -150 22 -149 24
rect -153 21 -149 22
rect -333 14 -332 16
rect -330 14 -329 16
rect -333 13 -329 14
rect -379 6 -378 8
rect -376 6 -375 8
rect -379 5 -375 6
rect -404 -10 -403 -8
rect -401 -10 -400 -8
rect -404 -11 -400 -10
rect -129 -8 -125 95
rect -129 -10 -128 -8
rect -126 -10 -125 -8
rect -129 -11 -125 -10
rect -119 56 -115 101
rect -104 100 -100 101
rect -104 98 -103 100
rect -101 98 -100 100
rect -104 64 -100 98
rect -104 62 -103 64
rect -101 62 -100 64
rect -104 61 -100 62
rect -119 54 -118 56
rect -116 54 -115 56
rect -119 -16 -115 54
rect -94 32 -90 101
rect -78 100 -74 101
rect -78 98 -77 100
rect -75 98 -74 100
rect -78 48 -74 98
rect -65 94 -61 95
rect -65 92 -64 94
rect -62 92 -61 94
rect -65 64 -61 92
rect -65 62 -64 64
rect -62 62 -61 64
rect -65 61 -61 62
rect -78 46 -77 48
rect -75 46 -74 48
rect -78 45 -74 46
rect -57 48 -53 109
rect -3 111 1 112
rect -3 109 -2 111
rect 0 109 1 111
rect 123 111 127 112
rect 123 109 124 111
rect 126 109 127 111
rect -24 101 -20 102
rect -24 99 -23 101
rect -21 99 -20 101
rect -57 46 -56 48
rect -54 46 -53 48
rect -57 45 -53 46
rect -48 96 -44 97
rect -48 94 -47 96
rect -45 94 -44 96
rect -94 30 -93 32
rect -91 30 -90 32
rect -94 8 -90 30
rect -48 24 -44 94
rect -24 40 -20 99
rect -11 94 -7 95
rect -11 92 -10 94
rect -8 92 -7 94
rect -11 56 -7 92
rect -11 54 -10 56
rect -8 54 -7 56
rect -11 53 -7 54
rect -3 48 1 109
rect 56 108 60 109
rect 56 106 57 108
rect 59 106 60 108
rect 30 101 34 102
rect 30 99 31 101
rect 33 99 34 101
rect -3 46 -2 48
rect 0 46 1 48
rect -3 45 1 46
rect 6 96 10 97
rect 6 94 7 96
rect 9 94 10 96
rect -24 38 -23 40
rect -21 38 -20 40
rect -24 37 -20 38
rect -48 22 -47 24
rect -45 22 -44 24
rect -48 16 -44 22
rect 6 24 10 94
rect 30 64 34 99
rect 30 62 31 64
rect 33 62 34 64
rect 30 61 34 62
rect 40 100 44 101
rect 40 98 41 100
rect 43 98 44 100
rect 40 64 44 98
rect 40 62 41 64
rect 43 62 44 64
rect 40 61 44 62
rect 56 56 60 106
rect 87 108 91 109
rect 87 106 88 108
rect 90 106 91 108
rect 75 100 79 101
rect 75 98 76 100
rect 78 98 79 100
rect 64 95 68 96
rect 64 93 65 95
rect 67 93 68 95
rect 64 64 68 93
rect 64 62 65 64
rect 67 62 68 64
rect 64 61 68 62
rect 75 64 79 98
rect 75 62 76 64
rect 78 62 79 64
rect 75 61 79 62
rect 87 64 91 106
rect 115 94 119 95
rect 87 62 88 64
rect 90 62 91 64
rect 56 54 57 56
rect 59 54 60 56
rect 56 53 60 54
rect 87 40 91 62
rect 99 93 103 94
rect 99 91 100 93
rect 102 91 103 93
rect 99 56 103 91
rect 99 54 100 56
rect 102 54 103 56
rect 99 53 103 54
rect 115 92 116 94
rect 118 92 119 94
rect 115 56 119 92
rect 115 54 116 56
rect 118 54 119 56
rect 115 53 119 54
rect 87 38 88 40
rect 90 38 91 40
rect 87 37 91 38
rect 123 32 127 109
rect 228 111 232 112
rect 228 109 229 111
rect 231 109 232 111
rect 123 30 124 32
rect 126 30 127 32
rect 123 29 127 30
rect 132 95 136 97
rect 132 93 133 95
rect 135 93 136 95
rect 6 22 7 24
rect 9 22 10 24
rect 6 21 10 22
rect 132 24 136 93
rect 142 70 146 104
rect 166 103 170 104
rect 166 101 167 103
rect 169 101 170 103
rect 191 103 195 105
rect 191 101 192 103
rect 194 101 195 103
rect 156 97 160 98
rect 156 95 157 97
rect 159 95 160 97
rect 156 40 160 95
rect 156 38 157 40
rect 159 38 160 40
rect 156 37 160 38
rect 166 56 170 101
rect 181 100 185 101
rect 181 98 182 100
rect 184 98 185 100
rect 181 64 185 98
rect 181 62 182 64
rect 184 62 185 64
rect 181 61 185 62
rect 166 54 167 56
rect 169 54 170 56
rect 132 22 133 24
rect 135 22 136 24
rect 132 21 136 22
rect -48 14 -47 16
rect -45 14 -44 16
rect -48 13 -44 14
rect -94 6 -93 8
rect -91 6 -90 8
rect -94 5 -90 6
rect 145 0 149 1
rect 145 -2 146 0
rect 148 -2 149 0
rect -119 -18 -118 -16
rect -116 -18 -115 -16
rect -119 -19 -115 -18
rect 136 -8 140 -7
rect 136 -10 137 -8
rect 139 -10 140 -8
rect -689 -26 -688 -24
rect -686 -26 -685 -24
rect -689 -27 -685 -26
rect 136 -24 140 -10
rect 145 -8 149 -2
rect 166 0 170 54
rect 191 32 195 101
rect 207 100 211 101
rect 207 98 208 100
rect 210 98 211 100
rect 207 48 211 98
rect 220 94 224 95
rect 220 92 221 94
rect 223 92 224 94
rect 220 64 224 92
rect 220 62 221 64
rect 223 62 224 64
rect 220 61 224 62
rect 207 46 208 48
rect 210 46 211 48
rect 207 45 211 46
rect 228 48 232 109
rect 282 111 286 112
rect 282 109 283 111
rect 285 109 286 111
rect 408 111 412 112
rect 408 109 409 111
rect 411 109 412 111
rect 261 101 265 102
rect 261 99 262 101
rect 264 99 265 101
rect 228 46 229 48
rect 231 46 232 48
rect 228 45 232 46
rect 237 96 241 97
rect 237 94 238 96
rect 240 94 241 96
rect 191 30 192 32
rect 194 30 195 32
rect 191 8 195 30
rect 191 6 192 8
rect 194 6 195 8
rect 191 5 195 6
rect 201 40 205 41
rect 201 38 202 40
rect 204 38 205 40
rect 201 8 205 38
rect 237 24 241 94
rect 261 40 265 99
rect 274 94 278 95
rect 274 92 275 94
rect 277 92 278 94
rect 274 56 278 92
rect 274 54 275 56
rect 277 54 278 56
rect 274 53 278 54
rect 282 48 286 109
rect 341 108 345 109
rect 341 106 342 108
rect 344 106 345 108
rect 315 101 319 102
rect 315 99 316 101
rect 318 99 319 101
rect 282 46 283 48
rect 285 46 286 48
rect 282 45 286 46
rect 291 96 295 97
rect 291 94 292 96
rect 294 94 295 96
rect 261 38 262 40
rect 264 38 265 40
rect 261 37 265 38
rect 237 22 238 24
rect 240 22 241 24
rect 237 16 241 22
rect 291 24 295 94
rect 315 64 319 99
rect 315 62 316 64
rect 318 62 319 64
rect 315 61 319 62
rect 325 100 329 101
rect 325 98 326 100
rect 328 98 329 100
rect 325 64 329 98
rect 325 62 326 64
rect 328 62 329 64
rect 325 61 329 62
rect 341 56 345 106
rect 372 108 376 109
rect 372 106 373 108
rect 375 106 376 108
rect 360 100 364 101
rect 360 98 361 100
rect 363 98 364 100
rect 349 95 353 96
rect 349 93 350 95
rect 352 93 353 95
rect 349 64 353 93
rect 349 62 350 64
rect 352 62 353 64
rect 349 61 353 62
rect 360 64 364 98
rect 360 62 361 64
rect 363 62 364 64
rect 360 61 364 62
rect 372 64 376 106
rect 400 94 404 95
rect 372 62 373 64
rect 375 62 376 64
rect 341 54 342 56
rect 344 54 345 56
rect 341 53 345 54
rect 372 40 376 62
rect 384 93 388 94
rect 384 91 385 93
rect 387 91 388 93
rect 384 56 388 91
rect 384 54 385 56
rect 387 54 388 56
rect 384 53 388 54
rect 400 92 401 94
rect 403 92 404 94
rect 400 56 404 92
rect 400 54 401 56
rect 403 54 404 56
rect 400 53 404 54
rect 372 38 373 40
rect 375 38 376 40
rect 372 37 376 38
rect 408 32 412 109
rect 488 111 492 112
rect 488 109 489 111
rect 491 109 492 111
rect 408 30 409 32
rect 411 30 412 32
rect 408 29 412 30
rect 417 95 421 97
rect 417 93 418 95
rect 420 93 421 95
rect 291 22 292 24
rect 294 22 295 24
rect 291 21 295 22
rect 417 24 421 93
rect 427 70 431 104
rect 454 101 458 102
rect 454 99 455 101
rect 457 99 458 101
rect 441 97 445 98
rect 441 95 442 97
rect 444 95 445 97
rect 417 22 418 24
rect 420 22 421 24
rect 417 21 421 22
rect 441 24 445 95
rect 441 22 442 24
rect 444 22 445 24
rect 441 21 445 22
rect 454 48 458 99
rect 454 46 455 48
rect 457 46 458 48
rect 237 14 238 16
rect 240 14 241 16
rect 237 13 241 14
rect 454 16 458 46
rect 478 94 482 95
rect 478 92 479 94
rect 481 92 482 94
rect 478 32 482 92
rect 488 56 492 109
rect 548 111 552 112
rect 548 109 549 111
rect 551 109 552 111
rect 514 101 518 102
rect 514 99 515 101
rect 517 99 518 101
rect 496 96 504 97
rect 496 94 497 96
rect 499 94 504 96
rect 496 93 504 94
rect 499 65 504 93
rect 499 64 503 65
rect 499 62 500 64
rect 502 62 503 64
rect 499 61 503 62
rect 488 54 489 56
rect 491 54 492 56
rect 488 53 492 54
rect 478 30 479 32
rect 481 30 482 32
rect 478 29 482 30
rect 514 48 518 99
rect 514 46 515 48
rect 517 46 518 48
rect 454 14 455 16
rect 457 14 458 16
rect 454 13 458 14
rect 201 6 202 8
rect 204 6 205 8
rect 201 5 205 6
rect 166 -2 167 0
rect 169 -2 170 0
rect 166 -3 170 -2
rect 145 -10 146 -8
rect 148 -10 149 -8
rect 145 -11 149 -10
rect 469 -8 473 -7
rect 469 -10 470 -8
rect 472 -10 473 -8
rect 136 -26 137 -24
rect 139 -26 140 -24
rect 136 -27 140 -26
rect -699 -114 -698 -112
rect -696 -114 -695 -112
rect -699 -302 -695 -114
rect -689 -40 -685 -39
rect -689 -42 -688 -40
rect -686 -42 -685 -40
rect -689 -120 -685 -42
rect 156 -40 160 -39
rect 156 -42 157 -40
rect 159 -42 160 -40
rect -119 -48 -115 -47
rect -119 -50 -118 -48
rect -116 -50 -115 -48
rect -404 -56 -400 -55
rect -404 -58 -403 -56
rect -401 -58 -400 -56
rect -414 -64 -410 -63
rect -414 -66 -413 -64
rect -411 -66 -410 -64
rect -689 -122 -688 -120
rect -686 -122 -685 -120
rect -689 -167 -685 -122
rect -664 -72 -660 -71
rect -664 -74 -663 -72
rect -661 -74 -660 -72
rect -664 -96 -660 -74
rect -664 -98 -663 -96
rect -661 -98 -660 -96
rect -664 -112 -660 -98
rect -618 -80 -614 -79
rect -618 -82 -617 -80
rect -615 -82 -614 -80
rect -618 -88 -614 -82
rect -618 -90 -617 -88
rect -615 -90 -614 -88
rect -664 -114 -663 -112
rect -661 -114 -660 -112
rect -674 -128 -670 -127
rect -674 -130 -673 -128
rect -671 -130 -670 -128
rect -674 -164 -670 -130
rect -674 -166 -673 -164
rect -671 -166 -670 -164
rect -674 -167 -670 -166
rect -664 -167 -660 -114
rect -648 -112 -644 -111
rect -648 -114 -647 -112
rect -645 -114 -644 -112
rect -648 -164 -644 -114
rect -627 -112 -623 -111
rect -627 -114 -626 -112
rect -624 -114 -623 -112
rect -635 -128 -631 -127
rect -635 -130 -634 -128
rect -632 -130 -631 -128
rect -635 -158 -631 -130
rect -635 -160 -634 -158
rect -632 -160 -631 -158
rect -635 -161 -631 -160
rect -648 -166 -647 -164
rect -645 -166 -644 -164
rect -648 -167 -644 -166
rect -689 -169 -688 -167
rect -686 -169 -685 -167
rect -689 -170 -685 -169
rect -664 -169 -663 -167
rect -661 -169 -660 -167
rect -664 -171 -660 -169
rect -627 -175 -623 -114
rect -618 -160 -614 -90
rect -564 -88 -560 -87
rect -564 -90 -563 -88
rect -561 -90 -560 -88
rect -618 -162 -617 -160
rect -615 -162 -614 -160
rect -618 -163 -614 -162
rect -594 -104 -590 -103
rect -594 -106 -593 -104
rect -591 -106 -590 -104
rect -594 -165 -590 -106
rect -573 -112 -569 -111
rect -573 -114 -572 -112
rect -570 -114 -569 -112
rect -581 -120 -577 -119
rect -581 -122 -580 -120
rect -578 -122 -577 -120
rect -581 -158 -577 -122
rect -581 -160 -580 -158
rect -578 -160 -577 -158
rect -581 -161 -577 -160
rect -594 -167 -593 -165
rect -591 -167 -590 -165
rect -594 -168 -590 -167
rect -627 -177 -626 -175
rect -624 -177 -623 -175
rect -627 -178 -623 -177
rect -573 -175 -569 -114
rect -564 -160 -560 -90
rect -438 -88 -434 -87
rect -438 -90 -437 -88
rect -435 -90 -434 -88
rect -447 -96 -443 -95
rect -447 -98 -446 -96
rect -444 -98 -443 -96
rect -483 -104 -479 -103
rect -483 -106 -482 -104
rect -480 -106 -479 -104
rect -514 -120 -510 -119
rect -514 -122 -513 -120
rect -511 -122 -510 -120
rect -564 -162 -563 -160
rect -561 -162 -560 -160
rect -564 -163 -560 -162
rect -540 -128 -536 -127
rect -540 -130 -539 -128
rect -537 -130 -536 -128
rect -540 -165 -536 -130
rect -540 -167 -539 -165
rect -537 -167 -536 -165
rect -530 -128 -526 -127
rect -530 -130 -529 -128
rect -527 -130 -526 -128
rect -530 -164 -526 -130
rect -530 -166 -529 -164
rect -527 -166 -526 -164
rect -530 -167 -526 -166
rect -540 -168 -536 -167
rect -514 -172 -510 -122
rect -506 -128 -502 -127
rect -506 -130 -505 -128
rect -503 -130 -502 -128
rect -506 -159 -502 -130
rect -506 -161 -505 -159
rect -503 -161 -502 -159
rect -506 -162 -502 -161
rect -495 -128 -491 -127
rect -495 -130 -494 -128
rect -492 -130 -491 -128
rect -495 -164 -491 -130
rect -495 -166 -494 -164
rect -492 -166 -491 -164
rect -495 -167 -491 -166
rect -483 -128 -479 -106
rect -483 -130 -482 -128
rect -480 -130 -479 -128
rect -514 -174 -513 -172
rect -511 -174 -510 -172
rect -514 -175 -510 -174
rect -483 -172 -479 -130
rect -471 -120 -467 -119
rect -471 -122 -470 -120
rect -468 -122 -467 -120
rect -471 -157 -467 -122
rect -471 -159 -470 -157
rect -468 -159 -467 -157
rect -471 -160 -467 -159
rect -455 -120 -451 -119
rect -455 -122 -454 -120
rect -452 -122 -451 -120
rect -455 -158 -451 -122
rect -455 -160 -454 -158
rect -452 -160 -451 -158
rect -455 -161 -451 -160
rect -483 -174 -482 -172
rect -480 -174 -479 -172
rect -483 -175 -479 -174
rect -447 -175 -443 -98
rect -438 -159 -434 -90
rect -438 -161 -437 -159
rect -435 -161 -434 -159
rect -438 -163 -434 -161
rect -428 -170 -424 -136
rect -414 -161 -410 -66
rect -414 -163 -413 -161
rect -411 -163 -410 -161
rect -414 -164 -410 -163
rect -404 -120 -400 -58
rect -129 -56 -125 -55
rect -129 -58 -128 -56
rect -126 -58 -125 -56
rect -404 -122 -403 -120
rect -401 -122 -400 -120
rect -404 -167 -400 -122
rect -379 -72 -375 -71
rect -379 -74 -378 -72
rect -376 -74 -375 -72
rect -379 -96 -375 -74
rect -379 -98 -378 -96
rect -376 -98 -375 -96
rect -389 -128 -385 -127
rect -389 -130 -388 -128
rect -386 -130 -385 -128
rect -389 -164 -385 -130
rect -389 -166 -388 -164
rect -386 -166 -385 -164
rect -389 -167 -385 -166
rect -379 -167 -375 -98
rect -333 -80 -329 -79
rect -333 -82 -332 -80
rect -330 -82 -329 -80
rect -333 -88 -329 -82
rect -333 -90 -332 -88
rect -330 -90 -329 -88
rect -363 -112 -359 -111
rect -363 -114 -362 -112
rect -360 -114 -359 -112
rect -363 -164 -359 -114
rect -342 -112 -338 -111
rect -342 -114 -341 -112
rect -339 -114 -338 -112
rect -350 -128 -346 -127
rect -350 -130 -349 -128
rect -347 -130 -346 -128
rect -350 -158 -346 -130
rect -350 -160 -349 -158
rect -347 -160 -346 -158
rect -350 -161 -346 -160
rect -363 -166 -362 -164
rect -360 -166 -359 -164
rect -363 -167 -359 -166
rect -404 -169 -403 -167
rect -401 -169 -400 -167
rect -404 -170 -400 -169
rect -379 -169 -378 -167
rect -376 -169 -375 -167
rect -379 -171 -375 -169
rect -573 -177 -572 -175
rect -570 -177 -569 -175
rect -573 -178 -569 -177
rect -447 -177 -446 -175
rect -444 -177 -443 -175
rect -447 -178 -443 -177
rect -342 -175 -338 -114
rect -333 -160 -329 -90
rect -279 -88 -275 -87
rect -279 -90 -278 -88
rect -276 -90 -275 -88
rect -333 -162 -332 -160
rect -330 -162 -329 -160
rect -333 -163 -329 -162
rect -309 -104 -305 -103
rect -309 -106 -308 -104
rect -306 -106 -305 -104
rect -309 -165 -305 -106
rect -288 -112 -284 -111
rect -288 -114 -287 -112
rect -285 -114 -284 -112
rect -296 -120 -292 -119
rect -296 -122 -295 -120
rect -293 -122 -292 -120
rect -296 -158 -292 -122
rect -296 -160 -295 -158
rect -293 -160 -292 -158
rect -296 -161 -292 -160
rect -309 -167 -308 -165
rect -306 -167 -305 -165
rect -309 -168 -305 -167
rect -342 -177 -341 -175
rect -339 -177 -338 -175
rect -342 -178 -338 -177
rect -288 -175 -284 -114
rect -279 -160 -275 -90
rect -153 -88 -149 -87
rect -153 -90 -152 -88
rect -150 -90 -149 -88
rect -162 -96 -158 -95
rect -162 -98 -161 -96
rect -159 -98 -158 -96
rect -198 -104 -194 -103
rect -198 -106 -197 -104
rect -195 -106 -194 -104
rect -229 -120 -225 -119
rect -229 -122 -228 -120
rect -226 -122 -225 -120
rect -279 -162 -278 -160
rect -276 -162 -275 -160
rect -279 -163 -275 -162
rect -255 -128 -251 -127
rect -255 -130 -254 -128
rect -252 -130 -251 -128
rect -255 -165 -251 -130
rect -255 -167 -254 -165
rect -252 -167 -251 -165
rect -245 -128 -241 -127
rect -245 -130 -244 -128
rect -242 -130 -241 -128
rect -245 -164 -241 -130
rect -245 -166 -244 -164
rect -242 -166 -241 -164
rect -245 -167 -241 -166
rect -255 -168 -251 -167
rect -229 -172 -225 -122
rect -221 -128 -217 -127
rect -221 -130 -220 -128
rect -218 -130 -217 -128
rect -221 -159 -217 -130
rect -221 -161 -220 -159
rect -218 -161 -217 -159
rect -221 -162 -217 -161
rect -210 -128 -206 -127
rect -210 -130 -209 -128
rect -207 -130 -206 -128
rect -210 -164 -206 -130
rect -210 -166 -209 -164
rect -207 -166 -206 -164
rect -210 -167 -206 -166
rect -198 -128 -194 -106
rect -198 -130 -197 -128
rect -195 -130 -194 -128
rect -229 -174 -228 -172
rect -226 -174 -225 -172
rect -229 -175 -225 -174
rect -198 -172 -194 -130
rect -186 -120 -182 -119
rect -186 -122 -185 -120
rect -183 -122 -182 -120
rect -186 -157 -182 -122
rect -186 -159 -185 -157
rect -183 -159 -182 -157
rect -186 -160 -182 -159
rect -170 -120 -166 -119
rect -170 -122 -169 -120
rect -167 -122 -166 -120
rect -170 -158 -166 -122
rect -170 -160 -169 -158
rect -167 -160 -166 -158
rect -170 -161 -166 -160
rect -198 -174 -197 -172
rect -195 -174 -194 -172
rect -198 -175 -194 -174
rect -162 -175 -158 -98
rect -153 -159 -149 -90
rect -153 -161 -152 -159
rect -150 -161 -149 -159
rect -153 -163 -149 -161
rect -143 -170 -139 -136
rect -129 -161 -125 -58
rect -129 -163 -128 -161
rect -126 -163 -125 -161
rect -129 -164 -125 -163
rect -119 -120 -115 -50
rect 140 -56 144 -55
rect 140 -58 141 -56
rect 143 -58 144 -56
rect -119 -122 -118 -120
rect -116 -122 -115 -120
rect -119 -167 -115 -122
rect -94 -72 -90 -71
rect -94 -74 -93 -72
rect -91 -74 -90 -72
rect -94 -96 -90 -74
rect -94 -98 -93 -96
rect -91 -98 -90 -96
rect -104 -128 -100 -127
rect -104 -130 -103 -128
rect -101 -130 -100 -128
rect -104 -164 -100 -130
rect -104 -166 -103 -164
rect -101 -166 -100 -164
rect -104 -167 -100 -166
rect -94 -167 -90 -98
rect -48 -80 -44 -79
rect -48 -82 -47 -80
rect -45 -82 -44 -80
rect -48 -88 -44 -82
rect -48 -90 -47 -88
rect -45 -90 -44 -88
rect -78 -112 -74 -111
rect -78 -114 -77 -112
rect -75 -114 -74 -112
rect -78 -164 -74 -114
rect -57 -112 -53 -111
rect -57 -114 -56 -112
rect -54 -114 -53 -112
rect -65 -128 -61 -127
rect -65 -130 -64 -128
rect -62 -130 -61 -128
rect -65 -158 -61 -130
rect -65 -160 -64 -158
rect -62 -160 -61 -158
rect -65 -161 -61 -160
rect -78 -166 -77 -164
rect -75 -166 -74 -164
rect -78 -167 -74 -166
rect -119 -169 -118 -167
rect -116 -169 -115 -167
rect -119 -170 -115 -169
rect -94 -169 -93 -167
rect -91 -169 -90 -167
rect -94 -171 -90 -169
rect -288 -177 -287 -175
rect -285 -177 -284 -175
rect -288 -178 -284 -177
rect -162 -177 -161 -175
rect -159 -177 -158 -175
rect -162 -178 -158 -177
rect -57 -175 -53 -114
rect -48 -160 -44 -90
rect 6 -88 10 -87
rect 6 -90 7 -88
rect 9 -90 10 -88
rect -48 -162 -47 -160
rect -45 -162 -44 -160
rect -48 -163 -44 -162
rect -24 -104 -20 -103
rect -24 -106 -23 -104
rect -21 -106 -20 -104
rect -24 -165 -20 -106
rect -3 -112 1 -111
rect -3 -114 -2 -112
rect 0 -114 1 -112
rect -11 -120 -7 -119
rect -11 -122 -10 -120
rect -8 -122 -7 -120
rect -11 -158 -7 -122
rect -11 -160 -10 -158
rect -8 -160 -7 -158
rect -11 -161 -7 -160
rect -24 -167 -23 -165
rect -21 -167 -20 -165
rect -24 -168 -20 -167
rect -57 -177 -56 -175
rect -54 -177 -53 -175
rect -57 -178 -53 -177
rect -3 -175 1 -114
rect 6 -160 10 -90
rect 132 -88 136 -87
rect 132 -90 133 -88
rect 135 -90 136 -88
rect 123 -96 127 -95
rect 123 -98 124 -96
rect 126 -98 127 -96
rect 87 -104 91 -103
rect 87 -106 88 -104
rect 90 -106 91 -104
rect 56 -120 60 -119
rect 56 -122 57 -120
rect 59 -122 60 -120
rect 6 -162 7 -160
rect 9 -162 10 -160
rect 6 -163 10 -162
rect 30 -128 34 -127
rect 30 -130 31 -128
rect 33 -130 34 -128
rect 30 -165 34 -130
rect 30 -167 31 -165
rect 33 -167 34 -165
rect 40 -128 44 -127
rect 40 -130 41 -128
rect 43 -130 44 -128
rect 40 -164 44 -130
rect 40 -166 41 -164
rect 43 -166 44 -164
rect 40 -167 44 -166
rect 30 -168 34 -167
rect 56 -172 60 -122
rect 64 -128 68 -127
rect 64 -130 65 -128
rect 67 -130 68 -128
rect 64 -159 68 -130
rect 64 -161 65 -159
rect 67 -161 68 -159
rect 64 -162 68 -161
rect 75 -128 79 -127
rect 75 -130 76 -128
rect 78 -130 79 -128
rect 75 -164 79 -130
rect 75 -166 76 -164
rect 78 -166 79 -164
rect 75 -167 79 -166
rect 87 -128 91 -106
rect 87 -130 88 -128
rect 90 -130 91 -128
rect 56 -174 57 -172
rect 59 -174 60 -172
rect 56 -175 60 -174
rect 87 -172 91 -130
rect 99 -120 103 -119
rect 99 -122 100 -120
rect 102 -122 103 -120
rect 99 -157 103 -122
rect 99 -159 100 -157
rect 102 -159 103 -157
rect 99 -160 103 -159
rect 115 -120 119 -119
rect 115 -122 116 -120
rect 118 -122 119 -120
rect 115 -158 119 -122
rect 115 -160 116 -158
rect 118 -160 119 -158
rect 115 -161 119 -160
rect 87 -174 88 -172
rect 90 -174 91 -172
rect 87 -175 91 -174
rect 123 -175 127 -98
rect 132 -159 136 -90
rect 140 -88 144 -58
rect 148 -56 152 -55
rect 148 -58 149 -56
rect 151 -58 152 -56
rect 148 -64 152 -58
rect 148 -66 149 -64
rect 151 -66 152 -64
rect 148 -67 152 -66
rect 140 -90 141 -88
rect 143 -90 144 -88
rect 140 -91 144 -90
rect 132 -161 133 -159
rect 135 -161 136 -159
rect 132 -163 136 -161
rect 142 -170 146 -136
rect 156 -161 160 -42
rect 459 -56 463 -55
rect 459 -58 460 -56
rect 462 -58 463 -56
rect 156 -163 157 -161
rect 159 -163 160 -161
rect 156 -164 160 -163
rect 166 -64 170 -63
rect 166 -66 167 -64
rect 169 -66 170 -64
rect 166 -120 170 -66
rect 166 -122 167 -120
rect 169 -122 170 -120
rect 166 -167 170 -122
rect 191 -72 195 -71
rect 191 -74 192 -72
rect 194 -74 195 -72
rect 191 -96 195 -74
rect 229 -72 233 -71
rect 229 -74 230 -72
rect 232 -74 233 -72
rect 229 -88 233 -74
rect 229 -90 230 -88
rect 232 -90 233 -88
rect 229 -91 233 -90
rect 237 -80 241 -79
rect 237 -82 238 -80
rect 240 -82 241 -80
rect 237 -88 241 -82
rect 237 -90 238 -88
rect 240 -90 241 -88
rect 191 -98 192 -96
rect 194 -98 195 -96
rect 181 -128 185 -127
rect 181 -130 182 -128
rect 184 -130 185 -128
rect 181 -164 185 -130
rect 181 -166 182 -164
rect 184 -166 185 -164
rect 181 -167 185 -166
rect 191 -167 195 -98
rect 207 -112 211 -111
rect 207 -114 208 -112
rect 210 -114 211 -112
rect 207 -164 211 -114
rect 228 -112 232 -111
rect 228 -114 229 -112
rect 231 -114 232 -112
rect 220 -128 224 -127
rect 220 -130 221 -128
rect 223 -130 224 -128
rect 220 -158 224 -130
rect 220 -160 221 -158
rect 223 -160 224 -158
rect 220 -161 224 -160
rect 207 -166 208 -164
rect 210 -166 211 -164
rect 207 -167 211 -166
rect 166 -169 167 -167
rect 169 -169 170 -167
rect 166 -170 170 -169
rect 191 -169 192 -167
rect 194 -169 195 -167
rect 191 -171 195 -169
rect -3 -177 -2 -175
rect 0 -177 1 -175
rect -3 -178 1 -177
rect 123 -177 124 -175
rect 126 -177 127 -175
rect 123 -178 127 -177
rect 228 -175 232 -114
rect 237 -160 241 -90
rect 291 -88 295 -87
rect 291 -90 292 -88
rect 294 -90 295 -88
rect 237 -162 238 -160
rect 240 -162 241 -160
rect 237 -163 241 -162
rect 261 -104 265 -103
rect 261 -106 262 -104
rect 264 -106 265 -104
rect 261 -165 265 -106
rect 282 -112 286 -111
rect 282 -114 283 -112
rect 285 -114 286 -112
rect 274 -120 278 -119
rect 274 -122 275 -120
rect 277 -122 278 -120
rect 274 -158 278 -122
rect 274 -160 275 -158
rect 277 -160 278 -158
rect 274 -161 278 -160
rect 261 -167 262 -165
rect 264 -167 265 -165
rect 261 -168 265 -167
rect 228 -177 229 -175
rect 231 -177 232 -175
rect 228 -178 232 -177
rect 282 -175 286 -114
rect 291 -160 295 -90
rect 417 -88 421 -87
rect 417 -90 418 -88
rect 420 -90 421 -88
rect 408 -96 412 -95
rect 408 -98 409 -96
rect 411 -98 412 -96
rect 372 -104 376 -103
rect 372 -106 373 -104
rect 375 -106 376 -104
rect 341 -120 345 -119
rect 341 -122 342 -120
rect 344 -122 345 -120
rect 291 -162 292 -160
rect 294 -162 295 -160
rect 291 -163 295 -162
rect 315 -128 319 -127
rect 315 -130 316 -128
rect 318 -130 319 -128
rect 315 -165 319 -130
rect 315 -167 316 -165
rect 318 -167 319 -165
rect 325 -128 329 -127
rect 325 -130 326 -128
rect 328 -130 329 -128
rect 325 -164 329 -130
rect 325 -166 326 -164
rect 328 -166 329 -164
rect 325 -167 329 -166
rect 315 -168 319 -167
rect 341 -172 345 -122
rect 349 -128 353 -127
rect 349 -130 350 -128
rect 352 -130 353 -128
rect 349 -159 353 -130
rect 349 -161 350 -159
rect 352 -161 353 -159
rect 349 -162 353 -161
rect 360 -128 364 -127
rect 360 -130 361 -128
rect 363 -130 364 -128
rect 360 -164 364 -130
rect 360 -166 361 -164
rect 363 -166 364 -164
rect 360 -167 364 -166
rect 372 -128 376 -106
rect 372 -130 373 -128
rect 375 -130 376 -128
rect 341 -174 342 -172
rect 344 -174 345 -172
rect 341 -175 345 -174
rect 372 -172 376 -130
rect 384 -120 388 -119
rect 384 -122 385 -120
rect 387 -122 388 -120
rect 384 -157 388 -122
rect 384 -159 385 -157
rect 387 -159 388 -157
rect 384 -160 388 -159
rect 400 -120 404 -119
rect 400 -122 401 -120
rect 403 -122 404 -120
rect 400 -158 404 -122
rect 400 -160 401 -158
rect 403 -160 404 -158
rect 400 -161 404 -160
rect 372 -174 373 -172
rect 375 -174 376 -172
rect 372 -175 376 -174
rect 408 -175 412 -98
rect 417 -159 421 -90
rect 441 -88 445 -87
rect 441 -90 442 -88
rect 444 -90 445 -88
rect 417 -161 418 -159
rect 420 -161 421 -159
rect 417 -163 421 -161
rect 427 -170 431 -136
rect 441 -161 445 -90
rect 441 -163 442 -161
rect 444 -163 445 -161
rect 441 -164 445 -163
rect 282 -177 283 -175
rect 285 -177 286 -175
rect 282 -178 286 -177
rect 408 -177 409 -175
rect 411 -177 412 -175
rect 408 -178 412 -177
rect 459 -179 463 -58
rect 469 -174 473 -10
rect 514 -80 518 46
rect 538 94 542 95
rect 538 92 539 94
rect 541 92 542 94
rect 538 40 542 92
rect 548 82 552 109
rect 564 97 568 172
rect 556 96 568 97
rect 556 94 557 96
rect 559 94 568 96
rect 556 93 568 94
rect 596 103 600 105
rect 596 101 597 103
rect 599 101 600 103
rect 548 78 555 82
rect 551 56 555 78
rect 559 78 564 93
rect 580 87 584 89
rect 580 85 581 87
rect 583 85 584 87
rect 559 64 563 78
rect 559 62 560 64
rect 562 62 563 64
rect 559 61 563 62
rect 551 54 552 56
rect 554 54 555 56
rect 551 53 555 54
rect 580 48 584 85
rect 596 56 600 101
rect 596 54 597 56
rect 599 54 600 56
rect 596 53 600 54
rect 580 46 581 48
rect 583 46 584 48
rect 580 45 584 46
rect 608 48 612 244
rect 624 238 628 239
rect 624 236 625 238
rect 627 236 628 238
rect 608 46 609 48
rect 611 46 612 48
rect 608 45 612 46
rect 616 230 620 231
rect 616 228 617 230
rect 619 228 620 230
rect 538 38 539 40
rect 541 38 542 40
rect 538 37 542 38
rect 616 40 620 228
rect 616 38 617 40
rect 619 38 620 40
rect 616 37 620 38
rect 624 32 628 236
rect 624 30 625 32
rect 627 30 628 32
rect 624 29 628 30
rect 514 -82 515 -80
rect 517 -82 518 -80
rect 514 -83 518 -82
rect 551 -24 555 -23
rect 551 -26 552 -24
rect 554 -26 555 -24
rect 498 -120 502 -119
rect 498 -122 499 -120
rect 501 -122 502 -120
rect 487 -128 491 -127
rect 487 -130 488 -128
rect 490 -130 491 -128
rect 487 -159 491 -130
rect 487 -161 488 -159
rect 490 -161 491 -159
rect 487 -162 491 -161
rect 469 -176 470 -174
rect 472 -176 473 -174
rect 469 -177 473 -176
rect 498 -175 502 -122
rect 534 -162 538 -161
rect 534 -164 535 -162
rect 537 -164 538 -162
rect 534 -165 538 -164
rect 498 -177 499 -175
rect 501 -177 502 -175
rect 498 -178 502 -177
rect 459 -181 460 -179
rect 462 -181 463 -179
rect 459 -182 463 -181
rect 551 -180 555 -26
rect 561 -72 565 -71
rect 561 -74 562 -72
rect 564 -74 565 -72
rect 561 -174 565 -74
rect 590 -104 594 -103
rect 590 -106 591 -104
rect 593 -106 594 -104
rect 579 -112 583 -111
rect 579 -114 580 -112
rect 582 -114 583 -112
rect 579 -159 583 -114
rect 579 -161 580 -159
rect 582 -161 583 -159
rect 579 -162 583 -161
rect 561 -176 562 -174
rect 564 -176 565 -174
rect 561 -177 565 -176
rect 590 -175 594 -106
rect 590 -177 591 -175
rect 593 -177 594 -175
rect 590 -178 594 -177
rect 551 -182 552 -180
rect 554 -182 555 -180
rect 551 -183 555 -182
rect 459 -235 463 -233
rect 459 -237 460 -235
rect 462 -237 463 -235
rect -627 -239 -623 -238
rect -627 -241 -626 -239
rect -624 -241 -623 -239
rect -699 -304 -698 -302
rect -696 -304 -695 -302
rect -699 -305 -695 -304
rect -689 -247 -685 -246
rect -689 -249 -688 -247
rect -686 -249 -685 -247
rect -664 -247 -660 -245
rect -664 -249 -663 -247
rect -661 -249 -660 -247
rect -689 -294 -685 -249
rect -674 -250 -670 -249
rect -674 -252 -673 -250
rect -671 -252 -670 -250
rect -674 -286 -670 -252
rect -674 -288 -673 -286
rect -671 -288 -670 -286
rect -674 -289 -670 -288
rect -689 -296 -688 -294
rect -686 -296 -685 -294
rect -707 -352 -706 -350
rect -704 -352 -703 -350
rect -707 -353 -703 -352
rect -715 -360 -714 -358
rect -712 -360 -711 -358
rect -715 -361 -711 -360
rect -689 -358 -685 -296
rect -664 -302 -660 -249
rect -664 -304 -663 -302
rect -661 -304 -660 -302
rect -664 -318 -660 -304
rect -648 -250 -644 -249
rect -648 -252 -647 -250
rect -645 -252 -644 -250
rect -648 -302 -644 -252
rect -635 -256 -631 -255
rect -635 -258 -634 -256
rect -632 -258 -631 -256
rect -635 -286 -631 -258
rect -635 -288 -634 -286
rect -632 -288 -631 -286
rect -635 -289 -631 -288
rect -648 -304 -647 -302
rect -645 -304 -644 -302
rect -648 -305 -644 -304
rect -627 -302 -623 -241
rect -573 -239 -569 -238
rect -573 -241 -572 -239
rect -570 -241 -569 -239
rect -447 -239 -443 -238
rect -447 -241 -446 -239
rect -444 -241 -443 -239
rect -594 -249 -590 -248
rect -594 -251 -593 -249
rect -591 -251 -590 -249
rect -627 -304 -626 -302
rect -624 -304 -623 -302
rect -627 -305 -623 -304
rect -618 -254 -614 -253
rect -618 -256 -617 -254
rect -615 -256 -614 -254
rect -664 -320 -663 -318
rect -661 -320 -660 -318
rect -664 -342 -660 -320
rect -618 -326 -614 -256
rect -594 -310 -590 -251
rect -581 -256 -577 -255
rect -581 -258 -580 -256
rect -578 -258 -577 -256
rect -581 -294 -577 -258
rect -581 -296 -580 -294
rect -578 -296 -577 -294
rect -581 -297 -577 -296
rect -573 -302 -569 -241
rect -514 -242 -510 -241
rect -514 -244 -513 -242
rect -511 -244 -510 -242
rect -540 -249 -536 -248
rect -540 -251 -539 -249
rect -537 -251 -536 -249
rect -573 -304 -572 -302
rect -570 -304 -569 -302
rect -573 -305 -569 -304
rect -564 -254 -560 -253
rect -564 -256 -563 -254
rect -561 -256 -560 -254
rect -594 -312 -593 -310
rect -591 -312 -590 -310
rect -594 -313 -590 -312
rect -618 -328 -617 -326
rect -615 -328 -614 -326
rect -618 -334 -614 -328
rect -564 -326 -560 -256
rect -540 -286 -536 -251
rect -540 -288 -539 -286
rect -537 -288 -536 -286
rect -540 -289 -536 -288
rect -530 -250 -526 -249
rect -530 -252 -529 -250
rect -527 -252 -526 -250
rect -530 -286 -526 -252
rect -530 -288 -529 -286
rect -527 -288 -526 -286
rect -530 -289 -526 -288
rect -514 -294 -510 -244
rect -483 -242 -479 -241
rect -483 -244 -482 -242
rect -480 -244 -479 -242
rect -495 -250 -491 -249
rect -495 -252 -494 -250
rect -492 -252 -491 -250
rect -506 -255 -502 -254
rect -506 -257 -505 -255
rect -503 -257 -502 -255
rect -506 -286 -502 -257
rect -506 -288 -505 -286
rect -503 -288 -502 -286
rect -506 -289 -502 -288
rect -495 -286 -491 -252
rect -495 -288 -494 -286
rect -492 -288 -491 -286
rect -495 -289 -491 -288
rect -483 -286 -479 -244
rect -455 -256 -451 -255
rect -483 -288 -482 -286
rect -480 -288 -479 -286
rect -514 -296 -513 -294
rect -511 -296 -510 -294
rect -514 -297 -510 -296
rect -483 -310 -479 -288
rect -471 -257 -467 -256
rect -471 -259 -470 -257
rect -468 -259 -467 -257
rect -471 -294 -467 -259
rect -471 -296 -470 -294
rect -468 -296 -467 -294
rect -471 -297 -467 -296
rect -455 -258 -454 -256
rect -452 -258 -451 -256
rect -455 -294 -451 -258
rect -455 -296 -454 -294
rect -452 -296 -451 -294
rect -455 -297 -451 -296
rect -483 -312 -482 -310
rect -480 -312 -479 -310
rect -483 -313 -479 -312
rect -447 -318 -443 -241
rect -342 -239 -338 -238
rect -342 -241 -341 -239
rect -339 -241 -338 -239
rect -447 -320 -446 -318
rect -444 -320 -443 -318
rect -447 -321 -443 -320
rect -438 -255 -434 -253
rect -438 -257 -437 -255
rect -435 -257 -434 -255
rect -564 -328 -563 -326
rect -561 -328 -560 -326
rect -564 -329 -560 -328
rect -438 -326 -434 -257
rect -428 -280 -424 -246
rect -404 -247 -400 -246
rect -404 -249 -403 -247
rect -401 -249 -400 -247
rect -379 -247 -375 -245
rect -379 -249 -378 -247
rect -376 -249 -375 -247
rect -414 -253 -410 -252
rect -414 -255 -413 -253
rect -411 -255 -410 -253
rect -438 -328 -437 -326
rect -435 -328 -434 -326
rect -438 -329 -434 -328
rect -618 -336 -617 -334
rect -615 -336 -614 -334
rect -618 -337 -614 -336
rect -664 -344 -663 -342
rect -661 -344 -660 -342
rect -664 -345 -660 -344
rect -689 -360 -688 -358
rect -686 -360 -685 -358
rect -689 -361 -685 -360
rect -414 -367 -410 -255
rect -404 -294 -400 -249
rect -389 -250 -385 -249
rect -389 -252 -388 -250
rect -386 -252 -385 -250
rect -389 -286 -385 -252
rect -389 -288 -388 -286
rect -386 -288 -385 -286
rect -389 -289 -385 -288
rect -404 -296 -403 -294
rect -401 -296 -400 -294
rect -404 -350 -400 -296
rect -379 -318 -375 -249
rect -363 -250 -359 -249
rect -363 -252 -362 -250
rect -360 -252 -359 -250
rect -363 -302 -359 -252
rect -350 -256 -346 -255
rect -350 -258 -349 -256
rect -347 -258 -346 -256
rect -350 -286 -346 -258
rect -350 -288 -349 -286
rect -347 -288 -346 -286
rect -350 -289 -346 -288
rect -363 -304 -362 -302
rect -360 -304 -359 -302
rect -363 -305 -359 -304
rect -342 -302 -338 -241
rect -288 -239 -284 -238
rect -288 -241 -287 -239
rect -285 -241 -284 -239
rect -162 -239 -158 -238
rect -162 -241 -161 -239
rect -159 -241 -158 -239
rect -309 -249 -305 -248
rect -309 -251 -308 -249
rect -306 -251 -305 -249
rect -342 -304 -341 -302
rect -339 -304 -338 -302
rect -342 -305 -338 -304
rect -333 -254 -329 -253
rect -333 -256 -332 -254
rect -330 -256 -329 -254
rect -379 -320 -378 -318
rect -376 -320 -375 -318
rect -379 -342 -375 -320
rect -333 -326 -329 -256
rect -309 -310 -305 -251
rect -296 -256 -292 -255
rect -296 -258 -295 -256
rect -293 -258 -292 -256
rect -296 -294 -292 -258
rect -296 -296 -295 -294
rect -293 -296 -292 -294
rect -296 -297 -292 -296
rect -288 -302 -284 -241
rect -229 -242 -225 -241
rect -229 -244 -228 -242
rect -226 -244 -225 -242
rect -255 -249 -251 -248
rect -255 -251 -254 -249
rect -252 -251 -251 -249
rect -288 -304 -287 -302
rect -285 -304 -284 -302
rect -288 -305 -284 -304
rect -279 -254 -275 -253
rect -279 -256 -278 -254
rect -276 -256 -275 -254
rect -309 -312 -308 -310
rect -306 -312 -305 -310
rect -309 -313 -305 -312
rect -333 -328 -332 -326
rect -330 -328 -329 -326
rect -333 -334 -329 -328
rect -279 -326 -275 -256
rect -255 -286 -251 -251
rect -255 -288 -254 -286
rect -252 -288 -251 -286
rect -255 -289 -251 -288
rect -245 -250 -241 -249
rect -245 -252 -244 -250
rect -242 -252 -241 -250
rect -245 -286 -241 -252
rect -245 -288 -244 -286
rect -242 -288 -241 -286
rect -245 -289 -241 -288
rect -229 -294 -225 -244
rect -198 -242 -194 -241
rect -198 -244 -197 -242
rect -195 -244 -194 -242
rect -210 -250 -206 -249
rect -210 -252 -209 -250
rect -207 -252 -206 -250
rect -221 -255 -217 -254
rect -221 -257 -220 -255
rect -218 -257 -217 -255
rect -221 -286 -217 -257
rect -221 -288 -220 -286
rect -218 -288 -217 -286
rect -221 -289 -217 -288
rect -210 -286 -206 -252
rect -210 -288 -209 -286
rect -207 -288 -206 -286
rect -210 -289 -206 -288
rect -198 -286 -194 -244
rect -170 -256 -166 -255
rect -198 -288 -197 -286
rect -195 -288 -194 -286
rect -229 -296 -228 -294
rect -226 -296 -225 -294
rect -229 -297 -225 -296
rect -198 -310 -194 -288
rect -186 -257 -182 -256
rect -186 -259 -185 -257
rect -183 -259 -182 -257
rect -186 -294 -182 -259
rect -186 -296 -185 -294
rect -183 -296 -182 -294
rect -186 -297 -182 -296
rect -170 -258 -169 -256
rect -167 -258 -166 -256
rect -170 -294 -166 -258
rect -170 -296 -169 -294
rect -167 -296 -166 -294
rect -170 -297 -166 -296
rect -198 -312 -197 -310
rect -195 -312 -194 -310
rect -198 -313 -194 -312
rect -162 -318 -158 -241
rect -57 -239 -53 -238
rect -57 -241 -56 -239
rect -54 -241 -53 -239
rect -162 -320 -161 -318
rect -159 -320 -158 -318
rect -162 -321 -158 -320
rect -153 -255 -149 -253
rect -153 -257 -152 -255
rect -150 -257 -149 -255
rect -279 -328 -278 -326
rect -276 -328 -275 -326
rect -279 -329 -275 -328
rect -153 -326 -149 -257
rect -143 -280 -139 -246
rect -119 -247 -115 -246
rect -119 -249 -118 -247
rect -116 -249 -115 -247
rect -94 -247 -90 -245
rect -94 -249 -93 -247
rect -91 -249 -90 -247
rect -129 -253 -125 -252
rect -129 -255 -128 -253
rect -126 -255 -125 -253
rect -153 -328 -152 -326
rect -150 -328 -149 -326
rect -153 -329 -149 -328
rect -333 -336 -332 -334
rect -330 -336 -329 -334
rect -333 -337 -329 -336
rect -379 -344 -378 -342
rect -376 -344 -375 -342
rect -379 -345 -375 -344
rect -404 -352 -403 -350
rect -401 -352 -400 -350
rect -404 -353 -400 -352
rect -129 -350 -125 -255
rect -129 -352 -128 -350
rect -126 -352 -125 -350
rect -129 -353 -125 -352
rect -119 -294 -115 -249
rect -104 -250 -100 -249
rect -104 -252 -103 -250
rect -101 -252 -100 -250
rect -104 -286 -100 -252
rect -104 -288 -103 -286
rect -101 -288 -100 -286
rect -104 -289 -100 -288
rect -119 -296 -118 -294
rect -116 -296 -115 -294
rect -119 -358 -115 -296
rect -94 -318 -90 -249
rect -78 -250 -74 -249
rect -78 -252 -77 -250
rect -75 -252 -74 -250
rect -78 -302 -74 -252
rect -65 -256 -61 -255
rect -65 -258 -64 -256
rect -62 -258 -61 -256
rect -65 -286 -61 -258
rect -65 -288 -64 -286
rect -62 -288 -61 -286
rect -65 -289 -61 -288
rect -78 -304 -77 -302
rect -75 -304 -74 -302
rect -78 -305 -74 -304
rect -57 -302 -53 -241
rect -3 -239 1 -238
rect -3 -241 -2 -239
rect 0 -241 1 -239
rect 123 -239 127 -238
rect 123 -241 124 -239
rect 126 -241 127 -239
rect -24 -249 -20 -248
rect -24 -251 -23 -249
rect -21 -251 -20 -249
rect -57 -304 -56 -302
rect -54 -304 -53 -302
rect -57 -305 -53 -304
rect -48 -254 -44 -253
rect -48 -256 -47 -254
rect -45 -256 -44 -254
rect -94 -320 -93 -318
rect -91 -320 -90 -318
rect -94 -342 -90 -320
rect -48 -326 -44 -256
rect -24 -310 -20 -251
rect -11 -256 -7 -255
rect -11 -258 -10 -256
rect -8 -258 -7 -256
rect -11 -294 -7 -258
rect -11 -296 -10 -294
rect -8 -296 -7 -294
rect -11 -297 -7 -296
rect -3 -302 1 -241
rect 56 -242 60 -241
rect 56 -244 57 -242
rect 59 -244 60 -242
rect 30 -249 34 -248
rect 30 -251 31 -249
rect 33 -251 34 -249
rect -3 -304 -2 -302
rect 0 -304 1 -302
rect -3 -305 1 -304
rect 6 -254 10 -253
rect 6 -256 7 -254
rect 9 -256 10 -254
rect -24 -312 -23 -310
rect -21 -312 -20 -310
rect -24 -313 -20 -312
rect -48 -328 -47 -326
rect -45 -328 -44 -326
rect -48 -334 -44 -328
rect 6 -326 10 -256
rect 30 -286 34 -251
rect 30 -288 31 -286
rect 33 -288 34 -286
rect 30 -289 34 -288
rect 40 -250 44 -249
rect 40 -252 41 -250
rect 43 -252 44 -250
rect 40 -286 44 -252
rect 40 -288 41 -286
rect 43 -288 44 -286
rect 40 -289 44 -288
rect 56 -294 60 -244
rect 87 -242 91 -241
rect 87 -244 88 -242
rect 90 -244 91 -242
rect 75 -250 79 -249
rect 75 -252 76 -250
rect 78 -252 79 -250
rect 64 -255 68 -254
rect 64 -257 65 -255
rect 67 -257 68 -255
rect 64 -286 68 -257
rect 64 -288 65 -286
rect 67 -288 68 -286
rect 64 -289 68 -288
rect 75 -286 79 -252
rect 75 -288 76 -286
rect 78 -288 79 -286
rect 75 -289 79 -288
rect 87 -286 91 -244
rect 115 -256 119 -255
rect 87 -288 88 -286
rect 90 -288 91 -286
rect 56 -296 57 -294
rect 59 -296 60 -294
rect 56 -297 60 -296
rect 87 -310 91 -288
rect 99 -257 103 -256
rect 99 -259 100 -257
rect 102 -259 103 -257
rect 99 -294 103 -259
rect 99 -296 100 -294
rect 102 -296 103 -294
rect 99 -297 103 -296
rect 115 -258 116 -256
rect 118 -258 119 -256
rect 115 -294 119 -258
rect 115 -296 116 -294
rect 118 -296 119 -294
rect 115 -297 119 -296
rect 87 -312 88 -310
rect 90 -312 91 -310
rect 87 -313 91 -312
rect 123 -318 127 -241
rect 228 -239 232 -238
rect 228 -241 229 -239
rect 231 -241 232 -239
rect 123 -320 124 -318
rect 126 -320 127 -318
rect 123 -321 127 -320
rect 132 -255 136 -253
rect 132 -257 133 -255
rect 135 -257 136 -255
rect 6 -328 7 -326
rect 9 -328 10 -326
rect 6 -329 10 -328
rect 132 -326 136 -257
rect 142 -280 146 -246
rect 166 -247 170 -246
rect 166 -249 167 -247
rect 169 -249 170 -247
rect 191 -247 195 -245
rect 191 -249 192 -247
rect 194 -249 195 -247
rect 156 -253 160 -252
rect 156 -255 157 -253
rect 159 -255 160 -253
rect 132 -328 133 -326
rect 135 -328 136 -326
rect 132 -329 136 -328
rect 156 -326 160 -255
rect 156 -328 157 -326
rect 159 -328 160 -326
rect 156 -329 160 -328
rect 166 -294 170 -249
rect 181 -250 185 -249
rect 181 -252 182 -250
rect 184 -252 185 -250
rect 181 -286 185 -252
rect 181 -288 182 -286
rect 184 -288 185 -286
rect 181 -289 185 -288
rect 166 -296 167 -294
rect 169 -296 170 -294
rect -48 -336 -47 -334
rect -45 -336 -44 -334
rect -48 -337 -44 -336
rect -94 -344 -93 -342
rect -91 -344 -90 -342
rect -94 -345 -90 -344
rect -119 -360 -118 -358
rect -116 -360 -115 -358
rect -119 -361 -115 -360
rect 157 -350 161 -349
rect 157 -352 158 -350
rect 160 -352 161 -350
rect -414 -369 -413 -367
rect -411 -369 -410 -367
rect -414 -370 -410 -369
rect 157 -375 161 -352
rect 166 -350 170 -296
rect 191 -318 195 -249
rect 207 -250 211 -249
rect 207 -252 208 -250
rect 210 -252 211 -250
rect 207 -302 211 -252
rect 220 -256 224 -255
rect 220 -258 221 -256
rect 223 -258 224 -256
rect 220 -286 224 -258
rect 220 -288 221 -286
rect 223 -288 224 -286
rect 220 -289 224 -288
rect 207 -304 208 -302
rect 210 -304 211 -302
rect 207 -305 211 -304
rect 228 -302 232 -241
rect 282 -239 286 -238
rect 282 -241 283 -239
rect 285 -241 286 -239
rect 408 -239 412 -238
rect 408 -241 409 -239
rect 411 -241 412 -239
rect 261 -249 265 -248
rect 261 -251 262 -249
rect 264 -251 265 -249
rect 228 -304 229 -302
rect 231 -304 232 -302
rect 228 -305 232 -304
rect 237 -254 241 -253
rect 237 -256 238 -254
rect 240 -256 241 -254
rect 191 -320 192 -318
rect 194 -320 195 -318
rect 191 -342 195 -320
rect 191 -344 192 -342
rect 194 -344 195 -342
rect 191 -345 195 -344
rect 199 -326 203 -325
rect 199 -328 200 -326
rect 202 -328 203 -326
rect 199 -342 203 -328
rect 237 -326 241 -256
rect 261 -310 265 -251
rect 274 -256 278 -255
rect 274 -258 275 -256
rect 277 -258 278 -256
rect 274 -294 278 -258
rect 274 -296 275 -294
rect 277 -296 278 -294
rect 274 -297 278 -296
rect 282 -302 286 -241
rect 341 -242 345 -241
rect 341 -244 342 -242
rect 344 -244 345 -242
rect 315 -249 319 -248
rect 315 -251 316 -249
rect 318 -251 319 -249
rect 282 -304 283 -302
rect 285 -304 286 -302
rect 282 -305 286 -304
rect 291 -254 295 -253
rect 291 -256 292 -254
rect 294 -256 295 -254
rect 261 -312 262 -310
rect 264 -312 265 -310
rect 261 -313 265 -312
rect 237 -328 238 -326
rect 240 -328 241 -326
rect 237 -334 241 -328
rect 291 -326 295 -256
rect 315 -286 319 -251
rect 315 -288 316 -286
rect 318 -288 319 -286
rect 315 -289 319 -288
rect 325 -250 329 -249
rect 325 -252 326 -250
rect 328 -252 329 -250
rect 325 -286 329 -252
rect 325 -288 326 -286
rect 328 -288 329 -286
rect 325 -289 329 -288
rect 341 -294 345 -244
rect 372 -242 376 -241
rect 372 -244 373 -242
rect 375 -244 376 -242
rect 360 -250 364 -249
rect 360 -252 361 -250
rect 363 -252 364 -250
rect 349 -255 353 -254
rect 349 -257 350 -255
rect 352 -257 353 -255
rect 349 -286 353 -257
rect 349 -288 350 -286
rect 352 -288 353 -286
rect 349 -289 353 -288
rect 360 -286 364 -252
rect 360 -288 361 -286
rect 363 -288 364 -286
rect 360 -289 364 -288
rect 372 -286 376 -244
rect 400 -256 404 -255
rect 372 -288 373 -286
rect 375 -288 376 -286
rect 341 -296 342 -294
rect 344 -296 345 -294
rect 341 -297 345 -296
rect 372 -310 376 -288
rect 384 -257 388 -256
rect 384 -259 385 -257
rect 387 -259 388 -257
rect 384 -294 388 -259
rect 384 -296 385 -294
rect 387 -296 388 -294
rect 384 -297 388 -296
rect 400 -258 401 -256
rect 403 -258 404 -256
rect 400 -294 404 -258
rect 400 -296 401 -294
rect 403 -296 404 -294
rect 400 -297 404 -296
rect 372 -312 373 -310
rect 375 -312 376 -310
rect 372 -313 376 -312
rect 408 -318 412 -241
rect 408 -320 409 -318
rect 411 -320 412 -318
rect 408 -321 412 -320
rect 417 -255 421 -253
rect 417 -257 418 -255
rect 420 -257 421 -255
rect 291 -328 292 -326
rect 294 -328 295 -326
rect 291 -329 295 -328
rect 417 -326 421 -257
rect 427 -280 431 -246
rect 441 -253 445 -252
rect 441 -255 442 -253
rect 444 -255 445 -253
rect 441 -295 445 -255
rect 459 -287 463 -237
rect 553 -235 557 -234
rect 553 -237 554 -235
rect 556 -237 557 -235
rect 459 -289 460 -287
rect 462 -289 463 -287
rect 459 -290 463 -289
rect 469 -240 473 -238
rect 469 -242 470 -240
rect 472 -242 473 -240
rect 441 -297 442 -295
rect 444 -297 445 -295
rect 441 -298 445 -297
rect 469 -303 473 -242
rect 492 -239 496 -238
rect 492 -241 493 -239
rect 495 -241 496 -239
rect 469 -305 470 -303
rect 472 -305 473 -303
rect 469 -306 473 -305
rect 481 -255 485 -254
rect 481 -257 482 -255
rect 484 -257 485 -255
rect 481 -311 485 -257
rect 481 -313 482 -311
rect 484 -313 485 -311
rect 481 -314 485 -313
rect 417 -328 418 -326
rect 420 -328 421 -326
rect 417 -329 421 -328
rect 237 -336 238 -334
rect 240 -336 241 -334
rect 237 -337 241 -336
rect 199 -344 200 -342
rect 202 -344 203 -342
rect 199 -345 203 -344
rect 492 -342 496 -241
rect 553 -295 557 -237
rect 553 -297 554 -295
rect 556 -297 557 -295
rect 553 -298 557 -297
rect 561 -241 565 -238
rect 561 -243 562 -241
rect 564 -243 565 -241
rect 561 -295 565 -243
rect 598 -239 602 -238
rect 598 -241 599 -239
rect 601 -241 602 -239
rect 561 -297 562 -295
rect 564 -297 565 -295
rect 561 -298 565 -297
rect 571 -255 575 -254
rect 571 -257 572 -255
rect 574 -257 575 -255
rect 571 -319 575 -257
rect 571 -321 572 -319
rect 574 -321 575 -319
rect 571 -322 575 -321
rect 598 -327 602 -241
rect 598 -329 599 -327
rect 601 -329 602 -327
rect 598 -330 602 -329
rect 632 -335 636 260
rect 632 -337 633 -335
rect 635 -337 636 -335
rect 632 -338 636 -337
rect 640 0 644 284
rect 640 -2 641 0
rect 643 -2 644 0
rect 640 -64 644 -2
rect 640 -66 641 -64
rect 643 -66 644 -64
rect 492 -344 493 -342
rect 495 -344 496 -342
rect 492 -345 496 -344
rect 166 -352 167 -350
rect 169 -352 170 -350
rect 166 -353 170 -352
rect 640 -350 644 -66
rect 640 -352 641 -350
rect 643 -352 644 -350
rect 640 -353 644 -352
rect 648 -16 652 292
rect 648 -18 649 -16
rect 651 -18 652 -16
rect 648 -48 652 -18
rect 648 -50 649 -48
rect 651 -50 652 -48
rect 648 -358 652 -50
rect 656 -128 660 300
rect 664 -104 668 308
rect 664 -106 665 -104
rect 667 -106 668 -104
rect 664 -107 668 -106
rect 672 -104 676 316
rect 680 278 684 279
rect 680 276 681 278
rect 683 276 684 278
rect 680 33 684 276
rect 737 211 744 214
rect 737 209 739 211
rect 741 209 744 211
rect 737 75 744 209
rect 737 73 740 75
rect 742 73 744 75
rect 680 31 681 33
rect 683 31 684 33
rect 680 30 684 31
rect 704 33 708 34
rect 704 31 705 33
rect 707 31 708 33
rect 680 8 684 9
rect 680 6 681 8
rect 683 6 684 8
rect 680 -96 684 6
rect 696 -40 700 -39
rect 696 -42 697 -40
rect 699 -42 700 -40
rect 680 -98 681 -96
rect 683 -98 684 -96
rect 680 -99 684 -98
rect 688 -96 692 -95
rect 688 -98 689 -96
rect 691 -98 692 -96
rect 672 -106 673 -104
rect 675 -106 676 -104
rect 672 -107 676 -106
rect 680 -104 684 -103
rect 680 -106 681 -104
rect 683 -106 684 -104
rect 672 -112 676 -111
rect 672 -114 673 -112
rect 675 -114 676 -112
rect 656 -130 657 -128
rect 659 -130 660 -128
rect 656 -131 660 -130
rect 664 -120 668 -119
rect 664 -122 665 -120
rect 667 -122 668 -120
rect 656 -150 660 -149
rect 656 -152 657 -150
rect 659 -152 660 -150
rect 656 -295 660 -152
rect 656 -297 657 -295
rect 659 -297 660 -295
rect 656 -298 660 -297
rect 648 -360 649 -358
rect 651 -360 652 -358
rect 648 -361 652 -360
rect 664 -367 668 -122
rect 664 -369 665 -367
rect 667 -369 668 -367
rect 664 -370 668 -369
rect 157 -377 158 -375
rect 160 -377 161 -375
rect 157 -378 161 -377
rect 672 -375 676 -114
rect 680 -287 684 -106
rect 680 -289 681 -287
rect 683 -289 684 -287
rect 680 -290 684 -289
rect 688 -303 692 -98
rect 688 -305 689 -303
rect 691 -305 692 -303
rect 688 -306 692 -305
rect 696 -311 700 -42
rect 704 -150 708 31
rect 720 24 724 25
rect 720 22 721 24
rect 723 22 724 24
rect 704 -152 705 -150
rect 707 -152 708 -150
rect 704 -153 708 -152
rect 712 -88 716 -87
rect 712 -90 713 -88
rect 715 -90 716 -88
rect 696 -313 697 -311
rect 699 -313 700 -311
rect 696 -314 700 -313
rect 704 -158 708 -157
rect 704 -160 705 -158
rect 707 -160 708 -158
rect 704 -319 708 -160
rect 712 -158 716 -90
rect 712 -160 713 -158
rect 715 -160 716 -158
rect 712 -161 716 -160
rect 704 -321 705 -319
rect 707 -321 708 -319
rect 704 -322 708 -321
rect 712 -166 716 -165
rect 712 -168 713 -166
rect 715 -168 716 -166
rect 712 -327 716 -168
rect 720 -166 724 22
rect 720 -168 721 -166
rect 723 -168 724 -166
rect 720 -169 724 -168
rect 737 -139 744 73
rect 737 -141 739 -139
rect 741 -141 744 -139
rect 737 -275 744 -141
rect 737 -277 739 -275
rect 741 -277 744 -275
rect 737 -280 744 -277
rect 712 -329 713 -327
rect 715 -329 716 -327
rect 712 -330 716 -329
rect 672 -377 673 -375
rect 675 -377 676 -375
rect 672 -378 676 -377
<< ptie >>
rect -689 209 -671 211
rect -689 207 -687 209
rect -685 207 -675 209
rect -673 207 -671 209
rect -689 205 -671 207
rect -663 209 -645 211
rect -663 207 -661 209
rect -659 207 -649 209
rect -647 207 -645 209
rect -663 205 -645 207
rect -597 209 -591 211
rect -597 207 -595 209
rect -593 207 -591 209
rect -597 205 -591 207
rect -543 209 -537 211
rect -543 207 -541 209
rect -539 207 -537 209
rect -543 205 -537 207
rect -529 209 -523 211
rect -529 207 -527 209
rect -525 207 -523 209
rect -529 205 -523 207
rect -494 209 -488 211
rect -494 207 -492 209
rect -490 207 -488 209
rect -494 205 -488 207
rect -417 209 -411 211
rect -417 207 -415 209
rect -413 207 -411 209
rect -417 205 -411 207
rect -404 209 -386 211
rect -404 207 -402 209
rect -400 207 -390 209
rect -388 207 -386 209
rect -404 205 -386 207
rect -378 209 -360 211
rect -378 207 -376 209
rect -374 207 -364 209
rect -362 207 -360 209
rect -378 205 -360 207
rect -312 209 -306 211
rect -312 207 -310 209
rect -308 207 -306 209
rect -312 205 -306 207
rect -258 209 -252 211
rect -258 207 -256 209
rect -254 207 -252 209
rect -258 205 -252 207
rect -244 209 -238 211
rect -244 207 -242 209
rect -240 207 -238 209
rect -244 205 -238 207
rect -209 209 -203 211
rect -209 207 -207 209
rect -205 207 -203 209
rect -209 205 -203 207
rect -132 209 -126 211
rect -132 207 -130 209
rect -128 207 -126 209
rect -132 205 -126 207
rect -119 209 -101 211
rect -119 207 -117 209
rect -115 207 -105 209
rect -103 207 -101 209
rect -119 205 -101 207
rect -93 209 -75 211
rect -93 207 -91 209
rect -89 207 -79 209
rect -77 207 -75 209
rect -93 205 -75 207
rect -27 209 -21 211
rect -27 207 -25 209
rect -23 207 -21 209
rect -27 205 -21 207
rect 27 209 33 211
rect 27 207 29 209
rect 31 207 33 209
rect 27 205 33 207
rect 41 209 47 211
rect 41 207 43 209
rect 45 207 47 209
rect 41 205 47 207
rect 76 209 82 211
rect 76 207 78 209
rect 80 207 82 209
rect 76 205 82 207
rect 153 209 159 211
rect 153 207 155 209
rect 157 207 159 209
rect 153 205 159 207
rect 166 209 184 211
rect 166 207 168 209
rect 170 207 180 209
rect 182 207 184 209
rect 166 205 184 207
rect 192 209 210 211
rect 192 207 194 209
rect 196 207 206 209
rect 208 207 210 209
rect 192 205 210 207
rect 258 209 264 211
rect 258 207 260 209
rect 262 207 264 209
rect 258 205 264 207
rect 312 209 318 211
rect 312 207 314 209
rect 316 207 318 209
rect 312 205 318 207
rect 326 209 332 211
rect 326 207 328 209
rect 330 207 332 209
rect 326 205 332 207
rect 361 209 367 211
rect 361 207 363 209
rect 365 207 367 209
rect 361 205 367 207
rect 438 209 444 211
rect 438 207 440 209
rect 442 207 444 209
rect 438 205 444 207
rect 455 209 461 211
rect 455 207 457 209
rect 459 207 461 209
rect 455 205 461 207
rect 515 209 521 211
rect 515 207 517 209
rect 519 207 521 209
rect 515 205 521 207
rect 581 209 599 211
rect 581 207 583 209
rect 585 207 595 209
rect 597 207 599 209
rect 581 205 599 207
rect -689 77 -671 79
rect -689 75 -687 77
rect -685 75 -675 77
rect -673 75 -671 77
rect -689 73 -671 75
rect -663 77 -645 79
rect -663 75 -661 77
rect -659 75 -649 77
rect -647 75 -645 77
rect -663 73 -645 75
rect -597 77 -591 79
rect -597 75 -595 77
rect -593 75 -591 77
rect -597 73 -591 75
rect -543 77 -537 79
rect -543 75 -541 77
rect -539 75 -537 77
rect -543 73 -537 75
rect -529 77 -523 79
rect -529 75 -527 77
rect -525 75 -523 77
rect -529 73 -523 75
rect -494 77 -488 79
rect -494 75 -492 77
rect -490 75 -488 77
rect -494 73 -488 75
rect -417 77 -411 79
rect -417 75 -415 77
rect -413 75 -411 77
rect -417 73 -411 75
rect -404 77 -386 79
rect -404 75 -402 77
rect -400 75 -390 77
rect -388 75 -386 77
rect -404 73 -386 75
rect -378 77 -360 79
rect -378 75 -376 77
rect -374 75 -364 77
rect -362 75 -360 77
rect -378 73 -360 75
rect -312 77 -306 79
rect -312 75 -310 77
rect -308 75 -306 77
rect -312 73 -306 75
rect -258 77 -252 79
rect -258 75 -256 77
rect -254 75 -252 77
rect -258 73 -252 75
rect -244 77 -238 79
rect -244 75 -242 77
rect -240 75 -238 77
rect -244 73 -238 75
rect -209 77 -203 79
rect -209 75 -207 77
rect -205 75 -203 77
rect -209 73 -203 75
rect -132 77 -126 79
rect -132 75 -130 77
rect -128 75 -126 77
rect -132 73 -126 75
rect -119 77 -101 79
rect -119 75 -117 77
rect -115 75 -105 77
rect -103 75 -101 77
rect -119 73 -101 75
rect -93 77 -75 79
rect -93 75 -91 77
rect -89 75 -79 77
rect -77 75 -75 77
rect -93 73 -75 75
rect -27 77 -21 79
rect -27 75 -25 77
rect -23 75 -21 77
rect -27 73 -21 75
rect 27 77 33 79
rect 27 75 29 77
rect 31 75 33 77
rect 27 73 33 75
rect 41 77 47 79
rect 41 75 43 77
rect 45 75 47 77
rect 41 73 47 75
rect 76 77 82 79
rect 76 75 78 77
rect 80 75 82 77
rect 76 73 82 75
rect 153 77 159 79
rect 153 75 155 77
rect 157 75 159 77
rect 153 73 159 75
rect 166 77 184 79
rect 166 75 168 77
rect 170 75 180 77
rect 182 75 184 77
rect 166 73 184 75
rect 192 77 210 79
rect 192 75 194 77
rect 196 75 206 77
rect 208 75 210 77
rect 192 73 210 75
rect 258 77 264 79
rect 258 75 260 77
rect 262 75 264 77
rect 258 73 264 75
rect 312 77 318 79
rect 312 75 314 77
rect 316 75 318 77
rect 312 73 318 75
rect 326 77 332 79
rect 326 75 328 77
rect 330 75 332 77
rect 326 73 332 75
rect 361 77 367 79
rect 361 75 363 77
rect 365 75 367 77
rect 361 73 367 75
rect 438 77 444 79
rect 438 75 440 77
rect 442 75 444 77
rect 438 73 444 75
rect 455 77 461 79
rect 455 75 457 77
rect 459 75 461 77
rect 455 73 461 75
rect 515 77 521 79
rect 515 75 517 77
rect 519 75 521 77
rect 515 73 521 75
rect 581 77 599 79
rect 581 75 583 77
rect 585 75 595 77
rect 597 75 599 77
rect 581 73 599 75
rect -689 -141 -671 -139
rect -689 -143 -687 -141
rect -685 -143 -675 -141
rect -673 -143 -671 -141
rect -689 -145 -671 -143
rect -663 -141 -645 -139
rect -663 -143 -661 -141
rect -659 -143 -649 -141
rect -647 -143 -645 -141
rect -663 -145 -645 -143
rect -597 -141 -591 -139
rect -597 -143 -595 -141
rect -593 -143 -591 -141
rect -597 -145 -591 -143
rect -543 -141 -537 -139
rect -543 -143 -541 -141
rect -539 -143 -537 -141
rect -543 -145 -537 -143
rect -529 -141 -523 -139
rect -529 -143 -527 -141
rect -525 -143 -523 -141
rect -529 -145 -523 -143
rect -494 -141 -488 -139
rect -494 -143 -492 -141
rect -490 -143 -488 -141
rect -494 -145 -488 -143
rect -417 -141 -411 -139
rect -417 -143 -415 -141
rect -413 -143 -411 -141
rect -417 -145 -411 -143
rect -404 -141 -386 -139
rect -404 -143 -402 -141
rect -400 -143 -390 -141
rect -388 -143 -386 -141
rect -404 -145 -386 -143
rect -378 -141 -360 -139
rect -378 -143 -376 -141
rect -374 -143 -364 -141
rect -362 -143 -360 -141
rect -378 -145 -360 -143
rect -312 -141 -306 -139
rect -312 -143 -310 -141
rect -308 -143 -306 -141
rect -312 -145 -306 -143
rect -258 -141 -252 -139
rect -258 -143 -256 -141
rect -254 -143 -252 -141
rect -258 -145 -252 -143
rect -244 -141 -238 -139
rect -244 -143 -242 -141
rect -240 -143 -238 -141
rect -244 -145 -238 -143
rect -209 -141 -203 -139
rect -209 -143 -207 -141
rect -205 -143 -203 -141
rect -209 -145 -203 -143
rect -132 -141 -126 -139
rect -132 -143 -130 -141
rect -128 -143 -126 -141
rect -132 -145 -126 -143
rect -119 -141 -101 -139
rect -119 -143 -117 -141
rect -115 -143 -105 -141
rect -103 -143 -101 -141
rect -119 -145 -101 -143
rect -93 -141 -75 -139
rect -93 -143 -91 -141
rect -89 -143 -79 -141
rect -77 -143 -75 -141
rect -93 -145 -75 -143
rect -27 -141 -21 -139
rect -27 -143 -25 -141
rect -23 -143 -21 -141
rect -27 -145 -21 -143
rect 27 -141 33 -139
rect 27 -143 29 -141
rect 31 -143 33 -141
rect 27 -145 33 -143
rect 41 -141 47 -139
rect 41 -143 43 -141
rect 45 -143 47 -141
rect 41 -145 47 -143
rect 76 -141 82 -139
rect 76 -143 78 -141
rect 80 -143 82 -141
rect 76 -145 82 -143
rect 153 -141 159 -139
rect 153 -143 155 -141
rect 157 -143 159 -141
rect 153 -145 159 -143
rect 166 -141 184 -139
rect 166 -143 168 -141
rect 170 -143 180 -141
rect 182 -143 184 -141
rect 166 -145 184 -143
rect 192 -141 210 -139
rect 192 -143 194 -141
rect 196 -143 206 -141
rect 208 -143 210 -141
rect 192 -145 210 -143
rect 258 -141 264 -139
rect 258 -143 260 -141
rect 262 -143 264 -141
rect 258 -145 264 -143
rect 312 -141 318 -139
rect 312 -143 314 -141
rect 316 -143 318 -141
rect 312 -145 318 -143
rect 326 -141 332 -139
rect 326 -143 328 -141
rect 330 -143 332 -141
rect 326 -145 332 -143
rect 361 -141 367 -139
rect 361 -143 363 -141
rect 365 -143 367 -141
rect 361 -145 367 -143
rect 438 -141 444 -139
rect 438 -143 440 -141
rect 442 -143 444 -141
rect 438 -145 444 -143
rect 459 -141 473 -139
rect 459 -143 461 -141
rect 463 -143 469 -141
rect 471 -143 473 -141
rect 459 -160 473 -143
rect 551 -141 565 -139
rect 551 -143 553 -141
rect 555 -143 561 -141
rect 563 -143 565 -141
rect 551 -160 565 -143
rect -689 -273 -671 -271
rect -689 -275 -687 -273
rect -685 -275 -675 -273
rect -673 -275 -671 -273
rect -689 -277 -671 -275
rect -663 -273 -645 -271
rect -663 -275 -661 -273
rect -659 -275 -649 -273
rect -647 -275 -645 -273
rect -663 -277 -645 -275
rect -597 -273 -591 -271
rect -597 -275 -595 -273
rect -593 -275 -591 -273
rect -597 -277 -591 -275
rect -543 -273 -537 -271
rect -543 -275 -541 -273
rect -539 -275 -537 -273
rect -543 -277 -537 -275
rect -529 -273 -523 -271
rect -529 -275 -527 -273
rect -525 -275 -523 -273
rect -529 -277 -523 -275
rect -494 -273 -488 -271
rect -494 -275 -492 -273
rect -490 -275 -488 -273
rect -494 -277 -488 -275
rect -417 -273 -411 -271
rect -417 -275 -415 -273
rect -413 -275 -411 -273
rect -417 -277 -411 -275
rect -404 -273 -386 -271
rect -404 -275 -402 -273
rect -400 -275 -390 -273
rect -388 -275 -386 -273
rect -404 -277 -386 -275
rect -378 -273 -360 -271
rect -378 -275 -376 -273
rect -374 -275 -364 -273
rect -362 -275 -360 -273
rect -378 -277 -360 -275
rect -312 -273 -306 -271
rect -312 -275 -310 -273
rect -308 -275 -306 -273
rect -312 -277 -306 -275
rect -258 -273 -252 -271
rect -258 -275 -256 -273
rect -254 -275 -252 -273
rect -258 -277 -252 -275
rect -244 -273 -238 -271
rect -244 -275 -242 -273
rect -240 -275 -238 -273
rect -244 -277 -238 -275
rect -209 -273 -203 -271
rect -209 -275 -207 -273
rect -205 -275 -203 -273
rect -209 -277 -203 -275
rect -132 -273 -126 -271
rect -132 -275 -130 -273
rect -128 -275 -126 -273
rect -132 -277 -126 -275
rect -119 -273 -101 -271
rect -119 -275 -117 -273
rect -115 -275 -105 -273
rect -103 -275 -101 -273
rect -119 -277 -101 -275
rect -93 -273 -75 -271
rect -93 -275 -91 -273
rect -89 -275 -79 -273
rect -77 -275 -75 -273
rect -93 -277 -75 -275
rect -27 -273 -21 -271
rect -27 -275 -25 -273
rect -23 -275 -21 -273
rect -27 -277 -21 -275
rect 27 -273 33 -271
rect 27 -275 29 -273
rect 31 -275 33 -273
rect 27 -277 33 -275
rect 41 -273 47 -271
rect 41 -275 43 -273
rect 45 -275 47 -273
rect 41 -277 47 -275
rect 76 -273 82 -271
rect 76 -275 78 -273
rect 80 -275 82 -273
rect 76 -277 82 -275
rect 153 -273 159 -271
rect 153 -275 155 -273
rect 157 -275 159 -273
rect 153 -277 159 -275
rect 166 -273 184 -271
rect 166 -275 168 -273
rect 170 -275 180 -273
rect 182 -275 184 -273
rect 166 -277 184 -275
rect 192 -273 210 -271
rect 192 -275 194 -273
rect 196 -275 206 -273
rect 208 -275 210 -273
rect 192 -277 210 -275
rect 258 -273 264 -271
rect 258 -275 260 -273
rect 262 -275 264 -273
rect 258 -277 264 -275
rect 312 -273 318 -271
rect 312 -275 314 -273
rect 316 -275 318 -273
rect 312 -277 318 -275
rect 326 -273 332 -271
rect 326 -275 328 -273
rect 330 -275 332 -273
rect 326 -277 332 -275
rect 361 -273 367 -271
rect 361 -275 363 -273
rect 365 -275 367 -273
rect 361 -277 367 -275
rect 438 -273 444 -271
rect 438 -275 440 -273
rect 442 -275 444 -273
rect 438 -277 444 -275
rect 459 -273 473 -256
rect 459 -275 461 -273
rect 463 -275 469 -273
rect 471 -275 473 -273
rect 459 -277 473 -275
rect 551 -273 565 -256
rect 551 -275 553 -273
rect 555 -275 561 -273
rect 563 -275 565 -273
rect 551 -277 565 -275
<< ntie >>
rect -689 149 -671 151
rect -689 147 -687 149
rect -685 147 -675 149
rect -673 147 -671 149
rect -689 145 -671 147
rect -663 149 -645 151
rect -663 147 -661 149
rect -659 147 -649 149
rect -647 147 -645 149
rect -663 145 -645 147
rect -641 149 -635 151
rect -641 147 -639 149
rect -637 147 -635 149
rect -641 145 -635 147
rect -587 149 -581 151
rect -587 147 -585 149
rect -583 147 -581 149
rect -587 145 -581 147
rect -461 149 -455 151
rect -461 147 -459 149
rect -457 147 -455 149
rect -461 145 -455 147
rect -404 149 -386 151
rect -404 147 -402 149
rect -400 147 -390 149
rect -388 147 -386 149
rect -404 145 -386 147
rect -378 149 -360 151
rect -378 147 -376 149
rect -374 147 -364 149
rect -362 147 -360 149
rect -378 145 -360 147
rect -356 149 -350 151
rect -356 147 -354 149
rect -352 147 -350 149
rect -356 145 -350 147
rect -302 149 -296 151
rect -302 147 -300 149
rect -298 147 -296 149
rect -302 145 -296 147
rect -176 149 -170 151
rect -176 147 -174 149
rect -172 147 -170 149
rect -176 145 -170 147
rect -119 149 -101 151
rect -119 147 -117 149
rect -115 147 -105 149
rect -103 147 -101 149
rect -119 145 -101 147
rect -93 149 -75 151
rect -93 147 -91 149
rect -89 147 -79 149
rect -77 147 -75 149
rect -93 145 -75 147
rect -71 149 -65 151
rect -71 147 -69 149
rect -67 147 -65 149
rect -71 145 -65 147
rect -17 149 -11 151
rect -17 147 -15 149
rect -13 147 -11 149
rect -17 145 -11 147
rect 109 149 115 151
rect 109 147 111 149
rect 113 147 115 149
rect 109 145 115 147
rect 166 149 184 151
rect 166 147 168 149
rect 170 147 180 149
rect 182 147 184 149
rect 166 145 184 147
rect 192 149 210 151
rect 192 147 194 149
rect 196 147 206 149
rect 208 147 210 149
rect 192 145 210 147
rect 214 149 220 151
rect 214 147 216 149
rect 218 147 220 149
rect 214 145 220 147
rect 268 149 274 151
rect 268 147 270 149
rect 272 147 274 149
rect 268 145 274 147
rect 394 149 400 151
rect 394 147 396 149
rect 398 147 400 149
rect 394 145 400 147
rect 499 149 505 151
rect 499 147 501 149
rect 503 147 505 149
rect 499 145 505 147
rect 559 149 565 151
rect 559 147 561 149
rect 563 147 565 149
rect 559 145 565 147
rect 581 149 599 151
rect 581 147 583 149
rect 585 147 595 149
rect 597 147 599 149
rect 581 145 599 147
rect -689 137 -671 139
rect -689 135 -687 137
rect -685 135 -675 137
rect -673 135 -671 137
rect -689 133 -671 135
rect -663 137 -645 139
rect -663 135 -661 137
rect -659 135 -649 137
rect -647 135 -645 137
rect -663 133 -645 135
rect -641 137 -635 139
rect -641 135 -639 137
rect -637 135 -635 137
rect -641 133 -635 135
rect -587 137 -581 139
rect -587 135 -585 137
rect -583 135 -581 137
rect -587 133 -581 135
rect -461 137 -455 139
rect -461 135 -459 137
rect -457 135 -455 137
rect -461 133 -455 135
rect -404 137 -386 139
rect -404 135 -402 137
rect -400 135 -390 137
rect -388 135 -386 137
rect -404 133 -386 135
rect -378 137 -360 139
rect -378 135 -376 137
rect -374 135 -364 137
rect -362 135 -360 137
rect -378 133 -360 135
rect -356 137 -350 139
rect -356 135 -354 137
rect -352 135 -350 137
rect -356 133 -350 135
rect -302 137 -296 139
rect -302 135 -300 137
rect -298 135 -296 137
rect -302 133 -296 135
rect -176 137 -170 139
rect -176 135 -174 137
rect -172 135 -170 137
rect -176 133 -170 135
rect -119 137 -101 139
rect -119 135 -117 137
rect -115 135 -105 137
rect -103 135 -101 137
rect -119 133 -101 135
rect -93 137 -75 139
rect -93 135 -91 137
rect -89 135 -79 137
rect -77 135 -75 137
rect -93 133 -75 135
rect -71 137 -65 139
rect -71 135 -69 137
rect -67 135 -65 137
rect -71 133 -65 135
rect -17 137 -11 139
rect -17 135 -15 137
rect -13 135 -11 137
rect -17 133 -11 135
rect 109 137 115 139
rect 109 135 111 137
rect 113 135 115 137
rect 109 133 115 135
rect 166 137 184 139
rect 166 135 168 137
rect 170 135 180 137
rect 182 135 184 137
rect 166 133 184 135
rect 192 137 210 139
rect 192 135 194 137
rect 196 135 206 137
rect 208 135 210 137
rect 192 133 210 135
rect 214 137 220 139
rect 214 135 216 137
rect 218 135 220 137
rect 214 133 220 135
rect 268 137 274 139
rect 268 135 270 137
rect 272 135 274 137
rect 268 133 274 135
rect 394 137 400 139
rect 394 135 396 137
rect 398 135 400 137
rect 394 133 400 135
rect 499 137 505 139
rect 499 135 501 137
rect 503 135 505 137
rect 499 133 505 135
rect 559 137 565 139
rect 559 135 561 137
rect 563 135 565 137
rect 559 133 565 135
rect 581 137 599 139
rect 581 135 583 137
rect 585 135 595 137
rect 597 135 599 137
rect 581 133 599 135
rect -689 -201 -671 -199
rect -689 -203 -687 -201
rect -685 -203 -675 -201
rect -673 -203 -671 -201
rect -689 -205 -671 -203
rect -663 -201 -645 -199
rect -663 -203 -661 -201
rect -659 -203 -649 -201
rect -647 -203 -645 -201
rect -663 -205 -645 -203
rect -641 -201 -635 -199
rect -641 -203 -639 -201
rect -637 -203 -635 -201
rect -641 -205 -635 -203
rect -587 -201 -581 -199
rect -587 -203 -585 -201
rect -583 -203 -581 -201
rect -587 -205 -581 -203
rect -461 -201 -455 -199
rect -461 -203 -459 -201
rect -457 -203 -455 -201
rect -461 -205 -455 -203
rect -404 -201 -386 -199
rect -404 -203 -402 -201
rect -400 -203 -390 -201
rect -388 -203 -386 -201
rect -404 -205 -386 -203
rect -378 -201 -360 -199
rect -378 -203 -376 -201
rect -374 -203 -364 -201
rect -362 -203 -360 -201
rect -378 -205 -360 -203
rect -356 -201 -350 -199
rect -356 -203 -354 -201
rect -352 -203 -350 -201
rect -356 -205 -350 -203
rect -302 -201 -296 -199
rect -302 -203 -300 -201
rect -298 -203 -296 -201
rect -302 -205 -296 -203
rect -176 -201 -170 -199
rect -176 -203 -174 -201
rect -172 -203 -170 -201
rect -176 -205 -170 -203
rect -119 -201 -101 -199
rect -119 -203 -117 -201
rect -115 -203 -105 -201
rect -103 -203 -101 -201
rect -119 -205 -101 -203
rect -93 -201 -75 -199
rect -93 -203 -91 -201
rect -89 -203 -79 -201
rect -77 -203 -75 -201
rect -93 -205 -75 -203
rect -71 -201 -65 -199
rect -71 -203 -69 -201
rect -67 -203 -65 -201
rect -71 -205 -65 -203
rect -17 -201 -11 -199
rect -17 -203 -15 -201
rect -13 -203 -11 -201
rect -17 -205 -11 -203
rect 109 -201 115 -199
rect 109 -203 111 -201
rect 113 -203 115 -201
rect 109 -205 115 -203
rect 166 -201 184 -199
rect 166 -203 168 -201
rect 170 -203 180 -201
rect 182 -203 184 -201
rect 166 -205 184 -203
rect 192 -201 210 -199
rect 192 -203 194 -201
rect 196 -203 206 -201
rect 208 -203 210 -201
rect 192 -205 210 -203
rect 214 -201 220 -199
rect 214 -203 216 -201
rect 218 -203 220 -201
rect 214 -205 220 -203
rect 268 -201 274 -199
rect 268 -203 270 -201
rect 272 -203 274 -201
rect 268 -205 274 -203
rect 394 -201 400 -199
rect 394 -203 396 -201
rect 398 -203 400 -201
rect 394 -205 400 -203
rect 531 -201 537 -199
rect 531 -203 533 -201
rect 535 -203 537 -201
rect 531 -205 537 -203
rect 623 -201 629 -199
rect 623 -203 625 -201
rect 627 -203 629 -201
rect 623 -205 629 -203
rect -689 -213 -671 -211
rect -689 -215 -687 -213
rect -685 -215 -675 -213
rect -673 -215 -671 -213
rect -689 -217 -671 -215
rect -663 -213 -645 -211
rect -663 -215 -661 -213
rect -659 -215 -649 -213
rect -647 -215 -645 -213
rect -663 -217 -645 -215
rect -641 -213 -635 -211
rect -641 -215 -639 -213
rect -637 -215 -635 -213
rect -641 -217 -635 -215
rect -587 -213 -581 -211
rect -587 -215 -585 -213
rect -583 -215 -581 -213
rect -587 -217 -581 -215
rect -461 -213 -455 -211
rect -461 -215 -459 -213
rect -457 -215 -455 -213
rect -461 -217 -455 -215
rect -404 -213 -386 -211
rect -404 -215 -402 -213
rect -400 -215 -390 -213
rect -388 -215 -386 -213
rect -404 -217 -386 -215
rect -378 -213 -360 -211
rect -378 -215 -376 -213
rect -374 -215 -364 -213
rect -362 -215 -360 -213
rect -378 -217 -360 -215
rect -356 -213 -350 -211
rect -356 -215 -354 -213
rect -352 -215 -350 -213
rect -356 -217 -350 -215
rect -302 -213 -296 -211
rect -302 -215 -300 -213
rect -298 -215 -296 -213
rect -302 -217 -296 -215
rect -176 -213 -170 -211
rect -176 -215 -174 -213
rect -172 -215 -170 -213
rect -176 -217 -170 -215
rect -119 -213 -101 -211
rect -119 -215 -117 -213
rect -115 -215 -105 -213
rect -103 -215 -101 -213
rect -119 -217 -101 -215
rect -93 -213 -75 -211
rect -93 -215 -91 -213
rect -89 -215 -79 -213
rect -77 -215 -75 -213
rect -93 -217 -75 -215
rect -71 -213 -65 -211
rect -71 -215 -69 -213
rect -67 -215 -65 -213
rect -71 -217 -65 -215
rect -17 -213 -11 -211
rect -17 -215 -15 -213
rect -13 -215 -11 -213
rect -17 -217 -11 -215
rect 109 -213 115 -211
rect 109 -215 111 -213
rect 113 -215 115 -213
rect 109 -217 115 -215
rect 166 -213 184 -211
rect 166 -215 168 -213
rect 170 -215 180 -213
rect 182 -215 184 -213
rect 166 -217 184 -215
rect 192 -213 210 -211
rect 192 -215 194 -213
rect 196 -215 206 -213
rect 208 -215 210 -213
rect 192 -217 210 -215
rect 214 -213 220 -211
rect 214 -215 216 -213
rect 218 -215 220 -213
rect 214 -217 220 -215
rect 268 -213 274 -211
rect 268 -215 270 -213
rect 272 -215 274 -213
rect 268 -217 274 -215
rect 394 -213 400 -211
rect 394 -215 396 -213
rect 398 -215 400 -213
rect 394 -217 400 -215
rect 531 -213 537 -211
rect 531 -215 533 -213
rect 535 -215 537 -213
rect 531 -217 537 -215
rect 623 -213 629 -211
rect 623 -215 625 -213
rect 627 -215 629 -213
rect 623 -217 629 -215
<< nmos >>
rect -679 188 -677 197
rect -653 188 -651 197
rect -626 189 -624 202
rect -619 189 -617 202
rect -612 189 -610 202
rect -599 189 -597 198
rect -572 189 -570 202
rect -565 189 -563 202
rect -558 189 -556 202
rect -545 189 -543 198
rect -523 191 -521 199
rect -512 194 -510 202
rect -488 191 -486 199
rect -477 194 -475 202
rect -446 189 -444 202
rect -439 189 -437 202
rect -432 189 -430 202
rect -419 189 -417 198
rect -394 188 -392 197
rect -368 188 -366 197
rect -341 189 -339 202
rect -334 189 -332 202
rect -327 189 -325 202
rect -314 189 -312 198
rect -287 189 -285 202
rect -280 189 -278 202
rect -273 189 -271 202
rect -260 189 -258 198
rect -238 191 -236 199
rect -227 194 -225 202
rect -203 191 -201 199
rect -192 194 -190 202
rect -161 189 -159 202
rect -154 189 -152 202
rect -147 189 -145 202
rect -134 189 -132 198
rect -109 188 -107 197
rect -83 188 -81 197
rect -56 189 -54 202
rect -49 189 -47 202
rect -42 189 -40 202
rect -29 189 -27 198
rect -2 189 0 202
rect 5 189 7 202
rect 12 189 14 202
rect 25 189 27 198
rect 47 191 49 199
rect 58 194 60 202
rect 82 191 84 199
rect 93 194 95 202
rect 124 189 126 202
rect 131 189 133 202
rect 138 189 140 202
rect 151 189 153 198
rect 176 188 178 197
rect 202 188 204 197
rect 229 189 231 202
rect 236 189 238 202
rect 243 189 245 202
rect 256 189 258 198
rect 283 189 285 202
rect 290 189 292 202
rect 297 189 299 202
rect 310 189 312 198
rect 332 191 334 199
rect 343 194 345 202
rect 367 191 369 199
rect 378 194 380 202
rect 409 189 411 202
rect 416 189 418 202
rect 423 189 425 202
rect 436 189 438 198
rect 461 189 463 198
rect 474 189 476 202
rect 481 189 483 202
rect 488 189 490 202
rect 521 189 523 198
rect 534 189 536 202
rect 541 189 543 202
rect 548 189 550 202
rect 587 188 589 197
rect -679 87 -677 96
rect -653 87 -651 96
rect -626 82 -624 95
rect -619 82 -617 95
rect -612 82 -610 95
rect -599 86 -597 95
rect -572 82 -570 95
rect -565 82 -563 95
rect -558 82 -556 95
rect -545 86 -543 95
rect -523 85 -521 93
rect -512 82 -510 90
rect -488 85 -486 93
rect -477 82 -475 90
rect -446 82 -444 95
rect -439 82 -437 95
rect -432 82 -430 95
rect -419 86 -417 95
rect -394 87 -392 96
rect -368 87 -366 96
rect -341 82 -339 95
rect -334 82 -332 95
rect -327 82 -325 95
rect -314 86 -312 95
rect -287 82 -285 95
rect -280 82 -278 95
rect -273 82 -271 95
rect -260 86 -258 95
rect -238 85 -236 93
rect -227 82 -225 90
rect -203 85 -201 93
rect -192 82 -190 90
rect -161 82 -159 95
rect -154 82 -152 95
rect -147 82 -145 95
rect -134 86 -132 95
rect -109 87 -107 96
rect -83 87 -81 96
rect -56 82 -54 95
rect -49 82 -47 95
rect -42 82 -40 95
rect -29 86 -27 95
rect -2 82 0 95
rect 5 82 7 95
rect 12 82 14 95
rect 25 86 27 95
rect 47 85 49 93
rect 58 82 60 90
rect 82 85 84 93
rect 93 82 95 90
rect 124 82 126 95
rect 131 82 133 95
rect 138 82 140 95
rect 151 86 153 95
rect 176 87 178 96
rect 202 87 204 96
rect 229 82 231 95
rect 236 82 238 95
rect 243 82 245 95
rect 256 86 258 95
rect 283 82 285 95
rect 290 82 292 95
rect 297 82 299 95
rect 310 86 312 95
rect 332 85 334 93
rect 343 82 345 90
rect 367 85 369 93
rect 378 82 380 90
rect 409 82 411 95
rect 416 82 418 95
rect 423 82 425 95
rect 436 86 438 95
rect 461 86 463 95
rect 474 82 476 95
rect 481 82 483 95
rect 488 82 490 95
rect 521 86 523 95
rect 534 82 536 95
rect 541 82 543 95
rect 548 82 550 95
rect 587 87 589 96
rect -679 -162 -677 -153
rect -653 -162 -651 -153
rect -626 -161 -624 -148
rect -619 -161 -617 -148
rect -612 -161 -610 -148
rect -599 -161 -597 -152
rect -572 -161 -570 -148
rect -565 -161 -563 -148
rect -558 -161 -556 -148
rect -545 -161 -543 -152
rect -523 -159 -521 -151
rect -512 -156 -510 -148
rect -488 -159 -486 -151
rect -477 -156 -475 -148
rect -446 -161 -444 -148
rect -439 -161 -437 -148
rect -432 -161 -430 -148
rect -419 -161 -417 -152
rect -394 -162 -392 -153
rect -368 -162 -366 -153
rect -341 -161 -339 -148
rect -334 -161 -332 -148
rect -327 -161 -325 -148
rect -314 -161 -312 -152
rect -287 -161 -285 -148
rect -280 -161 -278 -148
rect -273 -161 -271 -148
rect -260 -161 -258 -152
rect -238 -159 -236 -151
rect -227 -156 -225 -148
rect -203 -159 -201 -151
rect -192 -156 -190 -148
rect -161 -161 -159 -148
rect -154 -161 -152 -148
rect -147 -161 -145 -148
rect -134 -161 -132 -152
rect -109 -162 -107 -153
rect -83 -162 -81 -153
rect -56 -161 -54 -148
rect -49 -161 -47 -148
rect -42 -161 -40 -148
rect -29 -161 -27 -152
rect -2 -161 0 -148
rect 5 -161 7 -148
rect 12 -161 14 -148
rect 25 -161 27 -152
rect 47 -159 49 -151
rect 58 -156 60 -148
rect 82 -159 84 -151
rect 93 -156 95 -148
rect 124 -161 126 -148
rect 131 -161 133 -148
rect 138 -161 140 -148
rect 151 -161 153 -152
rect 176 -162 178 -153
rect 202 -162 204 -153
rect 229 -161 231 -148
rect 236 -161 238 -148
rect 243 -161 245 -148
rect 256 -161 258 -152
rect 283 -161 285 -148
rect 290 -161 292 -148
rect 297 -161 299 -148
rect 310 -161 312 -152
rect 332 -159 334 -151
rect 343 -156 345 -148
rect 367 -159 369 -151
rect 378 -156 380 -148
rect 409 -161 411 -148
rect 416 -161 418 -148
rect 423 -161 425 -148
rect 436 -161 438 -152
rect 485 -154 487 -148
rect 495 -154 497 -148
rect 507 -154 509 -148
rect 517 -154 519 -148
rect 529 -157 531 -148
rect 577 -154 579 -148
rect 587 -154 589 -148
rect 599 -154 601 -148
rect 609 -154 611 -148
rect 621 -157 623 -148
rect -679 -263 -677 -254
rect -653 -263 -651 -254
rect -626 -268 -624 -255
rect -619 -268 -617 -255
rect -612 -268 -610 -255
rect -599 -264 -597 -255
rect -572 -268 -570 -255
rect -565 -268 -563 -255
rect -558 -268 -556 -255
rect -545 -264 -543 -255
rect -523 -265 -521 -257
rect -512 -268 -510 -260
rect -488 -265 -486 -257
rect -477 -268 -475 -260
rect -446 -268 -444 -255
rect -439 -268 -437 -255
rect -432 -268 -430 -255
rect -419 -264 -417 -255
rect -394 -263 -392 -254
rect -368 -263 -366 -254
rect -341 -268 -339 -255
rect -334 -268 -332 -255
rect -327 -268 -325 -255
rect -314 -264 -312 -255
rect -287 -268 -285 -255
rect -280 -268 -278 -255
rect -273 -268 -271 -255
rect -260 -264 -258 -255
rect -238 -265 -236 -257
rect -227 -268 -225 -260
rect -203 -265 -201 -257
rect -192 -268 -190 -260
rect -161 -268 -159 -255
rect -154 -268 -152 -255
rect -147 -268 -145 -255
rect -134 -264 -132 -255
rect -109 -263 -107 -254
rect -83 -263 -81 -254
rect -56 -268 -54 -255
rect -49 -268 -47 -255
rect -42 -268 -40 -255
rect -29 -264 -27 -255
rect -2 -268 0 -255
rect 5 -268 7 -255
rect 12 -268 14 -255
rect 25 -264 27 -255
rect 47 -265 49 -257
rect 58 -268 60 -260
rect 82 -265 84 -257
rect 93 -268 95 -260
rect 124 -268 126 -255
rect 131 -268 133 -255
rect 138 -268 140 -255
rect 151 -264 153 -255
rect 176 -263 178 -254
rect 202 -263 204 -254
rect 229 -268 231 -255
rect 236 -268 238 -255
rect 243 -268 245 -255
rect 256 -264 258 -255
rect 283 -268 285 -255
rect 290 -268 292 -255
rect 297 -268 299 -255
rect 310 -264 312 -255
rect 332 -265 334 -257
rect 343 -268 345 -260
rect 367 -265 369 -257
rect 378 -268 380 -260
rect 409 -268 411 -255
rect 416 -268 418 -255
rect 423 -268 425 -255
rect 436 -264 438 -255
rect 485 -268 487 -262
rect 495 -268 497 -262
rect 507 -268 509 -262
rect 517 -268 519 -262
rect 529 -268 531 -259
rect 577 -268 579 -262
rect 587 -268 589 -262
rect 599 -268 601 -262
rect 609 -268 611 -262
rect 621 -268 623 -259
<< pmos >>
rect -679 158 -677 176
rect -653 158 -651 176
rect -631 157 -629 170
rect -619 156 -617 169
rect -609 156 -607 169
rect -599 156 -597 174
rect -577 157 -575 170
rect -565 156 -563 169
rect -555 156 -553 169
rect -545 156 -543 174
rect -521 148 -519 176
rect -514 148 -512 176
rect -486 148 -484 176
rect -479 148 -477 176
rect -451 157 -449 170
rect -439 156 -437 169
rect -429 156 -427 169
rect -419 156 -417 174
rect -394 158 -392 176
rect -368 158 -366 176
rect -346 157 -344 170
rect -334 156 -332 169
rect -324 156 -322 169
rect -314 156 -312 174
rect -292 157 -290 170
rect -280 156 -278 169
rect -270 156 -268 169
rect -260 156 -258 174
rect -236 148 -234 176
rect -229 148 -227 176
rect -201 148 -199 176
rect -194 148 -192 176
rect -166 157 -164 170
rect -154 156 -152 169
rect -144 156 -142 169
rect -134 156 -132 174
rect -109 158 -107 176
rect -83 158 -81 176
rect -61 157 -59 170
rect -49 156 -47 169
rect -39 156 -37 169
rect -29 156 -27 174
rect -7 157 -5 170
rect 5 156 7 169
rect 15 156 17 169
rect 25 156 27 174
rect 49 148 51 176
rect 56 148 58 176
rect 84 148 86 176
rect 91 148 93 176
rect 119 157 121 170
rect 131 156 133 169
rect 141 156 143 169
rect 151 156 153 174
rect 176 158 178 176
rect 202 158 204 176
rect 224 157 226 170
rect 236 156 238 169
rect 246 156 248 169
rect 256 156 258 174
rect 278 157 280 170
rect 290 156 292 169
rect 300 156 302 169
rect 310 156 312 174
rect 334 148 336 176
rect 341 148 343 176
rect 369 148 371 176
rect 376 148 378 176
rect 404 157 406 170
rect 416 156 418 169
rect 426 156 428 169
rect 436 156 438 174
rect 461 156 463 174
rect 471 156 473 169
rect 481 156 483 169
rect 493 157 495 170
rect 521 156 523 174
rect 531 156 533 169
rect 541 156 543 169
rect 553 157 555 170
rect 587 158 589 176
rect -679 108 -677 126
rect -653 108 -651 126
rect -631 114 -629 127
rect -619 115 -617 128
rect -609 115 -607 128
rect -599 110 -597 128
rect -577 114 -575 127
rect -565 115 -563 128
rect -555 115 -553 128
rect -545 110 -543 128
rect -521 108 -519 136
rect -514 108 -512 136
rect -486 108 -484 136
rect -479 108 -477 136
rect -451 114 -449 127
rect -439 115 -437 128
rect -429 115 -427 128
rect -419 110 -417 128
rect -394 108 -392 126
rect -368 108 -366 126
rect -346 114 -344 127
rect -334 115 -332 128
rect -324 115 -322 128
rect -314 110 -312 128
rect -292 114 -290 127
rect -280 115 -278 128
rect -270 115 -268 128
rect -260 110 -258 128
rect -236 108 -234 136
rect -229 108 -227 136
rect -201 108 -199 136
rect -194 108 -192 136
rect -166 114 -164 127
rect -154 115 -152 128
rect -144 115 -142 128
rect -134 110 -132 128
rect -109 108 -107 126
rect -83 108 -81 126
rect -61 114 -59 127
rect -49 115 -47 128
rect -39 115 -37 128
rect -29 110 -27 128
rect -7 114 -5 127
rect 5 115 7 128
rect 15 115 17 128
rect 25 110 27 128
rect 49 108 51 136
rect 56 108 58 136
rect 84 108 86 136
rect 91 108 93 136
rect 119 114 121 127
rect 131 115 133 128
rect 141 115 143 128
rect 151 110 153 128
rect 176 108 178 126
rect 202 108 204 126
rect 224 114 226 127
rect 236 115 238 128
rect 246 115 248 128
rect 256 110 258 128
rect 278 114 280 127
rect 290 115 292 128
rect 300 115 302 128
rect 310 110 312 128
rect 334 108 336 136
rect 341 108 343 136
rect 369 108 371 136
rect 376 108 378 136
rect 404 114 406 127
rect 416 115 418 128
rect 426 115 428 128
rect 436 110 438 128
rect 461 110 463 128
rect 471 115 473 128
rect 481 115 483 128
rect 493 114 495 127
rect 521 110 523 128
rect 531 115 533 128
rect 541 115 543 128
rect 553 114 555 127
rect 587 108 589 126
rect -679 -192 -677 -174
rect -653 -192 -651 -174
rect -631 -193 -629 -180
rect -619 -194 -617 -181
rect -609 -194 -607 -181
rect -599 -194 -597 -176
rect -577 -193 -575 -180
rect -565 -194 -563 -181
rect -555 -194 -553 -181
rect -545 -194 -543 -176
rect -521 -202 -519 -174
rect -514 -202 -512 -174
rect -486 -202 -484 -174
rect -479 -202 -477 -174
rect -451 -193 -449 -180
rect -439 -194 -437 -181
rect -429 -194 -427 -181
rect -419 -194 -417 -176
rect -394 -192 -392 -174
rect -368 -192 -366 -174
rect -346 -193 -344 -180
rect -334 -194 -332 -181
rect -324 -194 -322 -181
rect -314 -194 -312 -176
rect -292 -193 -290 -180
rect -280 -194 -278 -181
rect -270 -194 -268 -181
rect -260 -194 -258 -176
rect -236 -202 -234 -174
rect -229 -202 -227 -174
rect -201 -202 -199 -174
rect -194 -202 -192 -174
rect -166 -193 -164 -180
rect -154 -194 -152 -181
rect -144 -194 -142 -181
rect -134 -194 -132 -176
rect -109 -192 -107 -174
rect -83 -192 -81 -174
rect -61 -193 -59 -180
rect -49 -194 -47 -181
rect -39 -194 -37 -181
rect -29 -194 -27 -176
rect -7 -193 -5 -180
rect 5 -194 7 -181
rect 15 -194 17 -181
rect 25 -194 27 -176
rect 49 -202 51 -174
rect 56 -202 58 -174
rect 84 -202 86 -174
rect 91 -202 93 -174
rect 119 -193 121 -180
rect 131 -194 133 -181
rect 141 -194 143 -181
rect 151 -194 153 -176
rect 176 -192 178 -174
rect 202 -192 204 -174
rect 224 -193 226 -180
rect 236 -194 238 -181
rect 246 -194 248 -181
rect 256 -194 258 -176
rect 278 -193 280 -180
rect 290 -194 292 -181
rect 300 -194 302 -181
rect 310 -194 312 -176
rect 334 -202 336 -174
rect 341 -202 343 -174
rect 369 -202 371 -174
rect 376 -202 378 -174
rect 404 -193 406 -180
rect 416 -194 418 -181
rect 426 -194 428 -181
rect 436 -194 438 -176
rect 465 -200 467 -182
rect 472 -200 474 -182
rect 479 -200 481 -182
rect 486 -200 488 -182
rect 496 -200 498 -182
rect 503 -200 505 -182
rect 510 -200 512 -182
rect 517 -200 519 -182
rect 529 -192 531 -174
rect 557 -200 559 -182
rect 564 -200 566 -182
rect 571 -200 573 -182
rect 578 -200 580 -182
rect 588 -200 590 -182
rect 595 -200 597 -182
rect 602 -200 604 -182
rect 609 -200 611 -182
rect 621 -192 623 -174
rect -679 -242 -677 -224
rect -653 -242 -651 -224
rect -631 -236 -629 -223
rect -619 -235 -617 -222
rect -609 -235 -607 -222
rect -599 -240 -597 -222
rect -577 -236 -575 -223
rect -565 -235 -563 -222
rect -555 -235 -553 -222
rect -545 -240 -543 -222
rect -521 -242 -519 -214
rect -514 -242 -512 -214
rect -486 -242 -484 -214
rect -479 -242 -477 -214
rect -451 -236 -449 -223
rect -439 -235 -437 -222
rect -429 -235 -427 -222
rect -419 -240 -417 -222
rect -394 -242 -392 -224
rect -368 -242 -366 -224
rect -346 -236 -344 -223
rect -334 -235 -332 -222
rect -324 -235 -322 -222
rect -314 -240 -312 -222
rect -292 -236 -290 -223
rect -280 -235 -278 -222
rect -270 -235 -268 -222
rect -260 -240 -258 -222
rect -236 -242 -234 -214
rect -229 -242 -227 -214
rect -201 -242 -199 -214
rect -194 -242 -192 -214
rect -166 -236 -164 -223
rect -154 -235 -152 -222
rect -144 -235 -142 -222
rect -134 -240 -132 -222
rect -109 -242 -107 -224
rect -83 -242 -81 -224
rect -61 -236 -59 -223
rect -49 -235 -47 -222
rect -39 -235 -37 -222
rect -29 -240 -27 -222
rect -7 -236 -5 -223
rect 5 -235 7 -222
rect 15 -235 17 -222
rect 25 -240 27 -222
rect 49 -242 51 -214
rect 56 -242 58 -214
rect 84 -242 86 -214
rect 91 -242 93 -214
rect 119 -236 121 -223
rect 131 -235 133 -222
rect 141 -235 143 -222
rect 151 -240 153 -222
rect 176 -242 178 -224
rect 202 -242 204 -224
rect 224 -236 226 -223
rect 236 -235 238 -222
rect 246 -235 248 -222
rect 256 -240 258 -222
rect 278 -236 280 -223
rect 290 -235 292 -222
rect 300 -235 302 -222
rect 310 -240 312 -222
rect 334 -242 336 -214
rect 341 -242 343 -214
rect 369 -242 371 -214
rect 376 -242 378 -214
rect 404 -236 406 -223
rect 416 -235 418 -222
rect 426 -235 428 -222
rect 436 -240 438 -222
rect 465 -234 467 -216
rect 472 -234 474 -216
rect 479 -234 481 -216
rect 486 -234 488 -216
rect 496 -234 498 -216
rect 503 -234 505 -216
rect 510 -234 512 -216
rect 517 -234 519 -216
rect 529 -242 531 -224
rect 557 -234 559 -216
rect 564 -234 566 -216
rect 571 -234 573 -216
rect 578 -234 580 -216
rect 588 -234 590 -216
rect 595 -234 597 -216
rect 602 -234 604 -216
rect 609 -234 611 -216
rect 621 -242 623 -224
<< polyct0 >>
rect -601 181 -599 183
rect -547 181 -545 183
rect -421 181 -419 183
rect -316 181 -314 183
rect -262 181 -260 183
rect -136 181 -134 183
rect -31 181 -29 183
rect 23 181 25 183
rect 149 181 151 183
rect 254 181 256 183
rect 308 181 310 183
rect 434 181 436 183
rect 463 181 465 183
rect 523 181 525 183
rect -601 101 -599 103
rect -547 101 -545 103
rect -421 101 -419 103
rect -316 101 -314 103
rect -262 101 -260 103
rect -136 101 -134 103
rect -31 101 -29 103
rect 23 101 25 103
rect 149 101 151 103
rect 254 101 256 103
rect 308 101 310 103
rect 434 101 436 103
rect 463 101 465 103
rect 523 101 525 103
rect -601 -169 -599 -167
rect -547 -169 -545 -167
rect -421 -169 -419 -167
rect -316 -169 -314 -167
rect -262 -169 -260 -167
rect -136 -169 -134 -167
rect -31 -169 -29 -167
rect 23 -169 25 -167
rect 149 -169 151 -167
rect 254 -169 256 -167
rect 308 -169 310 -167
rect 434 -169 436 -167
rect 527 -164 529 -162
rect 619 -164 621 -162
rect -601 -249 -599 -247
rect -547 -249 -545 -247
rect -421 -249 -419 -247
rect -316 -249 -314 -247
rect -262 -249 -260 -247
rect -136 -249 -134 -247
rect -31 -249 -29 -247
rect 23 -249 25 -247
rect 149 -249 151 -247
rect 254 -249 256 -247
rect 308 -249 310 -247
rect 434 -249 436 -247
rect 527 -254 529 -252
rect 619 -254 621 -252
<< polyct1 >>
rect -681 181 -679 183
rect -655 181 -653 183
rect -633 181 -631 183
rect -611 181 -609 183
rect -579 181 -577 183
rect -621 174 -619 176
rect -557 181 -555 183
rect -523 184 -521 186
rect -567 174 -565 176
rect -513 181 -511 183
rect -488 184 -486 186
rect -478 181 -476 183
rect -453 181 -451 183
rect -431 181 -429 183
rect -396 181 -394 183
rect -370 181 -368 183
rect -348 181 -346 183
rect -441 174 -439 176
rect -326 181 -324 183
rect -294 181 -292 183
rect -336 174 -334 176
rect -272 181 -270 183
rect -238 184 -236 186
rect -282 174 -280 176
rect -228 181 -226 183
rect -203 184 -201 186
rect -193 181 -191 183
rect -168 181 -166 183
rect -146 181 -144 183
rect -111 181 -109 183
rect -85 181 -83 183
rect -63 181 -61 183
rect -156 174 -154 176
rect -41 181 -39 183
rect -9 181 -7 183
rect -51 174 -49 176
rect 13 181 15 183
rect 47 184 49 186
rect 3 174 5 176
rect 57 181 59 183
rect 82 184 84 186
rect 92 181 94 183
rect 117 181 119 183
rect 139 181 141 183
rect 174 181 176 183
rect 200 181 202 183
rect 222 181 224 183
rect 129 174 131 176
rect 244 181 246 183
rect 276 181 278 183
rect 234 174 236 176
rect 298 181 300 183
rect 332 184 334 186
rect 288 174 290 176
rect 342 181 344 183
rect 367 184 369 186
rect 377 181 379 183
rect 402 181 404 183
rect 424 181 426 183
rect 414 174 416 176
rect 473 181 475 183
rect 495 181 497 183
rect 533 181 535 183
rect 483 174 485 176
rect 555 181 557 183
rect 589 181 591 183
rect 543 174 545 176
rect -621 108 -619 110
rect -681 101 -679 103
rect -655 101 -653 103
rect -633 101 -631 103
rect -567 108 -565 110
rect -611 101 -609 103
rect -579 101 -577 103
rect -557 101 -555 103
rect -523 98 -521 100
rect -513 101 -511 103
rect -441 108 -439 110
rect -488 98 -486 100
rect -478 101 -476 103
rect -453 101 -451 103
rect -336 108 -334 110
rect -431 101 -429 103
rect -396 101 -394 103
rect -370 101 -368 103
rect -348 101 -346 103
rect -282 108 -280 110
rect -326 101 -324 103
rect -294 101 -292 103
rect -272 101 -270 103
rect -238 98 -236 100
rect -228 101 -226 103
rect -156 108 -154 110
rect -203 98 -201 100
rect -193 101 -191 103
rect -168 101 -166 103
rect -51 108 -49 110
rect -146 101 -144 103
rect -111 101 -109 103
rect -85 101 -83 103
rect -63 101 -61 103
rect 3 108 5 110
rect -41 101 -39 103
rect -9 101 -7 103
rect 13 101 15 103
rect 47 98 49 100
rect 57 101 59 103
rect 129 108 131 110
rect 82 98 84 100
rect 92 101 94 103
rect 117 101 119 103
rect 234 108 236 110
rect 139 101 141 103
rect 174 101 176 103
rect 200 101 202 103
rect 222 101 224 103
rect 288 108 290 110
rect 244 101 246 103
rect 276 101 278 103
rect 298 101 300 103
rect 332 98 334 100
rect 342 101 344 103
rect 414 108 416 110
rect 367 98 369 100
rect 377 101 379 103
rect 402 101 404 103
rect 424 101 426 103
rect 483 108 485 110
rect 473 101 475 103
rect 543 108 545 110
rect 495 101 497 103
rect 533 101 535 103
rect 555 101 557 103
rect 589 101 591 103
rect -681 -169 -679 -167
rect -655 -169 -653 -167
rect -633 -169 -631 -167
rect -611 -169 -609 -167
rect -579 -169 -577 -167
rect -621 -176 -619 -174
rect -557 -169 -555 -167
rect -523 -166 -521 -164
rect -567 -176 -565 -174
rect -513 -169 -511 -167
rect -488 -166 -486 -164
rect -478 -169 -476 -167
rect -453 -169 -451 -167
rect -431 -169 -429 -167
rect -396 -169 -394 -167
rect -370 -169 -368 -167
rect -348 -169 -346 -167
rect -441 -176 -439 -174
rect -326 -169 -324 -167
rect -294 -169 -292 -167
rect -336 -176 -334 -174
rect -272 -169 -270 -167
rect -238 -166 -236 -164
rect -282 -176 -280 -174
rect -228 -169 -226 -167
rect -203 -166 -201 -164
rect -193 -169 -191 -167
rect -168 -169 -166 -167
rect -146 -169 -144 -167
rect -111 -169 -109 -167
rect -85 -169 -83 -167
rect -63 -169 -61 -167
rect -156 -176 -154 -174
rect -41 -169 -39 -167
rect -9 -169 -7 -167
rect -51 -176 -49 -174
rect 13 -169 15 -167
rect 47 -166 49 -164
rect 3 -176 5 -174
rect 57 -169 59 -167
rect 82 -166 84 -164
rect 92 -169 94 -167
rect 117 -169 119 -167
rect 139 -169 141 -167
rect 174 -169 176 -167
rect 200 -169 202 -167
rect 222 -169 224 -167
rect 129 -176 131 -174
rect 244 -169 246 -167
rect 276 -169 278 -167
rect 234 -176 236 -174
rect 298 -169 300 -167
rect 332 -166 334 -164
rect 288 -176 290 -174
rect 342 -169 344 -167
rect 367 -166 369 -164
rect 477 -161 479 -159
rect 377 -169 379 -167
rect 402 -169 404 -167
rect 424 -169 426 -167
rect 414 -176 416 -174
rect 471 -171 473 -169
rect 461 -177 463 -175
rect 493 -161 495 -159
rect 503 -165 505 -163
rect 487 -177 489 -175
rect 569 -161 571 -159
rect 518 -175 520 -173
rect 563 -171 565 -169
rect 553 -177 555 -175
rect 585 -161 587 -159
rect 595 -165 597 -163
rect 579 -177 581 -175
rect 610 -175 612 -173
rect -621 -242 -619 -240
rect -681 -249 -679 -247
rect -655 -249 -653 -247
rect -633 -249 -631 -247
rect -567 -242 -565 -240
rect -611 -249 -609 -247
rect -579 -249 -577 -247
rect -557 -249 -555 -247
rect -523 -252 -521 -250
rect -513 -249 -511 -247
rect -441 -242 -439 -240
rect -488 -252 -486 -250
rect -478 -249 -476 -247
rect -453 -249 -451 -247
rect -336 -242 -334 -240
rect -431 -249 -429 -247
rect -396 -249 -394 -247
rect -370 -249 -368 -247
rect -348 -249 -346 -247
rect -282 -242 -280 -240
rect -326 -249 -324 -247
rect -294 -249 -292 -247
rect -272 -249 -270 -247
rect -238 -252 -236 -250
rect -228 -249 -226 -247
rect -156 -242 -154 -240
rect -203 -252 -201 -250
rect -193 -249 -191 -247
rect -168 -249 -166 -247
rect -51 -242 -49 -240
rect -146 -249 -144 -247
rect -111 -249 -109 -247
rect -85 -249 -83 -247
rect -63 -249 -61 -247
rect 3 -242 5 -240
rect -41 -249 -39 -247
rect -9 -249 -7 -247
rect 13 -249 15 -247
rect 47 -252 49 -250
rect 57 -249 59 -247
rect 129 -242 131 -240
rect 82 -252 84 -250
rect 92 -249 94 -247
rect 117 -249 119 -247
rect 234 -242 236 -240
rect 139 -249 141 -247
rect 174 -249 176 -247
rect 200 -249 202 -247
rect 222 -249 224 -247
rect 288 -242 290 -240
rect 244 -249 246 -247
rect 276 -249 278 -247
rect 298 -249 300 -247
rect 332 -252 334 -250
rect 342 -249 344 -247
rect 414 -242 416 -240
rect 367 -252 369 -250
rect 377 -249 379 -247
rect 402 -249 404 -247
rect 461 -241 463 -239
rect 424 -249 426 -247
rect 471 -247 473 -245
rect 477 -257 479 -255
rect 487 -241 489 -239
rect 518 -243 520 -241
rect 553 -241 555 -239
rect 503 -253 505 -251
rect 493 -257 495 -255
rect 563 -247 565 -245
rect 569 -257 571 -255
rect 579 -241 581 -239
rect 610 -243 612 -241
rect 595 -253 597 -251
rect 585 -257 587 -255
<< ndifct0 >>
rect -631 198 -629 200
rect -688 193 -686 195
rect -662 193 -660 195
rect -577 198 -575 200
rect -528 195 -526 197
rect -493 195 -491 197
rect -451 198 -449 200
rect -346 198 -344 200
rect -403 193 -401 195
rect -377 193 -375 195
rect -292 198 -290 200
rect -243 195 -241 197
rect -208 195 -206 197
rect -166 198 -164 200
rect -61 198 -59 200
rect -118 193 -116 195
rect -92 193 -90 195
rect -7 198 -5 200
rect 42 195 44 197
rect 77 195 79 197
rect 119 198 121 200
rect 224 198 226 200
rect 167 193 169 195
rect 193 193 195 195
rect 278 198 280 200
rect 327 195 329 197
rect 362 195 364 197
rect 404 198 406 200
rect 493 198 495 200
rect 553 198 555 200
rect 596 193 598 195
rect -688 89 -686 91
rect -662 89 -660 91
rect -631 84 -629 86
rect -577 84 -575 86
rect -528 87 -526 89
rect -493 87 -491 89
rect -451 84 -449 86
rect -403 89 -401 91
rect -377 89 -375 91
rect -346 84 -344 86
rect -292 84 -290 86
rect -243 87 -241 89
rect -208 87 -206 89
rect -166 84 -164 86
rect -118 89 -116 91
rect -92 89 -90 91
rect -61 84 -59 86
rect -7 84 -5 86
rect 42 87 44 89
rect 77 87 79 89
rect 119 84 121 86
rect 167 89 169 91
rect 193 89 195 91
rect 224 84 226 86
rect 278 84 280 86
rect 327 87 329 89
rect 362 87 364 89
rect 404 84 406 86
rect 493 84 495 86
rect 596 89 598 91
rect 553 84 555 86
rect -631 -152 -629 -150
rect -688 -157 -686 -155
rect -662 -157 -660 -155
rect -577 -152 -575 -150
rect -528 -155 -526 -153
rect -493 -155 -491 -153
rect -451 -152 -449 -150
rect -346 -152 -344 -150
rect -403 -157 -401 -155
rect -377 -157 -375 -155
rect -292 -152 -290 -150
rect -243 -155 -241 -153
rect -208 -155 -206 -153
rect -166 -152 -164 -150
rect -61 -152 -59 -150
rect -118 -157 -116 -155
rect -92 -157 -90 -155
rect -7 -152 -5 -150
rect 42 -155 44 -153
rect 77 -155 79 -153
rect 119 -152 121 -150
rect 224 -152 226 -150
rect 167 -157 169 -155
rect 193 -157 195 -155
rect 278 -152 280 -150
rect 327 -155 329 -153
rect 362 -155 364 -153
rect 404 -152 406 -150
rect 490 -152 492 -150
rect 512 -152 514 -150
rect 582 -152 584 -150
rect 604 -152 606 -150
rect -688 -261 -686 -259
rect -662 -261 -660 -259
rect -631 -266 -629 -264
rect -577 -266 -575 -264
rect -528 -263 -526 -261
rect -493 -263 -491 -261
rect -451 -266 -449 -264
rect -403 -261 -401 -259
rect -377 -261 -375 -259
rect -346 -266 -344 -264
rect -292 -266 -290 -264
rect -243 -263 -241 -261
rect -208 -263 -206 -261
rect -166 -266 -164 -264
rect -118 -261 -116 -259
rect -92 -261 -90 -259
rect -61 -266 -59 -264
rect -7 -266 -5 -264
rect 42 -263 44 -261
rect 77 -263 79 -261
rect 119 -266 121 -264
rect 167 -261 169 -259
rect 193 -261 195 -259
rect 224 -266 226 -264
rect 278 -266 280 -264
rect 327 -263 329 -261
rect 362 -263 364 -261
rect 404 -266 406 -264
rect 490 -266 492 -264
rect 512 -266 514 -264
rect 582 -266 584 -264
rect 604 -266 606 -264
<< ndifct1 >>
rect -605 207 -603 209
rect -551 207 -549 209
rect -674 190 -672 192
rect -648 190 -646 192
rect -506 207 -504 209
rect -594 191 -592 193
rect -471 207 -469 209
rect -425 207 -423 209
rect -540 191 -538 193
rect -517 198 -515 200
rect -320 207 -318 209
rect -482 198 -480 200
rect -266 207 -264 209
rect -414 191 -412 193
rect -389 190 -387 192
rect -363 190 -361 192
rect -221 207 -219 209
rect -309 191 -307 193
rect -186 207 -184 209
rect -140 207 -138 209
rect -255 191 -253 193
rect -232 198 -230 200
rect -35 207 -33 209
rect -197 198 -195 200
rect 19 207 21 209
rect -129 191 -127 193
rect -104 190 -102 192
rect -78 190 -76 192
rect 64 207 66 209
rect -24 191 -22 193
rect 99 207 101 209
rect 145 207 147 209
rect 30 191 32 193
rect 53 198 55 200
rect 250 207 252 209
rect 88 198 90 200
rect 304 207 306 209
rect 156 191 158 193
rect 181 190 183 192
rect 207 190 209 192
rect 349 207 351 209
rect 261 191 263 193
rect 384 207 386 209
rect 430 207 432 209
rect 315 191 317 193
rect 338 198 340 200
rect 467 207 469 209
rect 373 198 375 200
rect 527 207 529 209
rect 441 191 443 193
rect 456 191 458 193
rect 516 191 518 193
rect 582 190 584 192
rect -674 92 -672 94
rect -648 92 -646 94
rect -594 91 -592 93
rect -540 91 -538 93
rect -605 75 -603 77
rect -517 84 -515 86
rect -551 75 -549 77
rect -482 84 -480 86
rect -414 91 -412 93
rect -389 92 -387 94
rect -363 92 -361 94
rect -506 75 -504 77
rect -309 91 -307 93
rect -471 75 -469 77
rect -425 75 -423 77
rect -255 91 -253 93
rect -320 75 -318 77
rect -232 84 -230 86
rect -266 75 -264 77
rect -197 84 -195 86
rect -129 91 -127 93
rect -104 92 -102 94
rect -78 92 -76 94
rect -221 75 -219 77
rect -24 91 -22 93
rect -186 75 -184 77
rect -140 75 -138 77
rect 30 91 32 93
rect -35 75 -33 77
rect 53 84 55 86
rect 19 75 21 77
rect 88 84 90 86
rect 156 91 158 93
rect 181 92 183 94
rect 207 92 209 94
rect 64 75 66 77
rect 261 91 263 93
rect 99 75 101 77
rect 145 75 147 77
rect 315 91 317 93
rect 250 75 252 77
rect 338 84 340 86
rect 304 75 306 77
rect 373 84 375 86
rect 441 91 443 93
rect 456 91 458 93
rect 349 75 351 77
rect 516 91 518 93
rect 384 75 386 77
rect 430 75 432 77
rect 582 92 584 94
rect 467 75 469 77
rect 527 75 529 77
rect -605 -143 -603 -141
rect -551 -143 -549 -141
rect -674 -160 -672 -158
rect -648 -160 -646 -158
rect -506 -143 -504 -141
rect -594 -159 -592 -157
rect -471 -143 -469 -141
rect -425 -143 -423 -141
rect -540 -159 -538 -157
rect -517 -152 -515 -150
rect -320 -143 -318 -141
rect -482 -152 -480 -150
rect -266 -143 -264 -141
rect -414 -159 -412 -157
rect -389 -160 -387 -158
rect -363 -160 -361 -158
rect -221 -143 -219 -141
rect -309 -159 -307 -157
rect -186 -143 -184 -141
rect -140 -143 -138 -141
rect -255 -159 -253 -157
rect -232 -152 -230 -150
rect -35 -143 -33 -141
rect -197 -152 -195 -150
rect 19 -143 21 -141
rect -129 -159 -127 -157
rect -104 -160 -102 -158
rect -78 -160 -76 -158
rect 64 -143 66 -141
rect -24 -159 -22 -157
rect 99 -143 101 -141
rect 145 -143 147 -141
rect 30 -159 32 -157
rect 53 -152 55 -150
rect 250 -143 252 -141
rect 88 -152 90 -150
rect 304 -143 306 -141
rect 156 -159 158 -157
rect 181 -160 183 -158
rect 207 -160 209 -158
rect 349 -143 351 -141
rect 261 -159 263 -157
rect 384 -143 386 -141
rect 430 -143 432 -141
rect 315 -159 317 -157
rect 338 -152 340 -150
rect 373 -152 375 -150
rect 441 -159 443 -157
rect 479 -143 481 -141
rect 501 -143 503 -141
rect 523 -143 525 -141
rect 534 -152 536 -150
rect 571 -143 573 -141
rect 593 -143 595 -141
rect 615 -143 617 -141
rect 626 -152 628 -150
rect -674 -258 -672 -256
rect -648 -258 -646 -256
rect -594 -259 -592 -257
rect -540 -259 -538 -257
rect -605 -275 -603 -273
rect -517 -266 -515 -264
rect -551 -275 -549 -273
rect -482 -266 -480 -264
rect -414 -259 -412 -257
rect -389 -258 -387 -256
rect -363 -258 -361 -256
rect -506 -275 -504 -273
rect -309 -259 -307 -257
rect -471 -275 -469 -273
rect -425 -275 -423 -273
rect -255 -259 -253 -257
rect -320 -275 -318 -273
rect -232 -266 -230 -264
rect -266 -275 -264 -273
rect -197 -266 -195 -264
rect -129 -259 -127 -257
rect -104 -258 -102 -256
rect -78 -258 -76 -256
rect -221 -275 -219 -273
rect -24 -259 -22 -257
rect -186 -275 -184 -273
rect -140 -275 -138 -273
rect 30 -259 32 -257
rect -35 -275 -33 -273
rect 53 -266 55 -264
rect 19 -275 21 -273
rect 88 -266 90 -264
rect 156 -259 158 -257
rect 181 -258 183 -256
rect 207 -258 209 -256
rect 64 -275 66 -273
rect 261 -259 263 -257
rect 99 -275 101 -273
rect 145 -275 147 -273
rect 315 -259 317 -257
rect 250 -275 252 -273
rect 338 -266 340 -264
rect 304 -275 306 -273
rect 373 -266 375 -264
rect 441 -259 443 -257
rect 349 -275 351 -273
rect 384 -275 386 -273
rect 430 -275 432 -273
rect 534 -266 536 -264
rect 479 -275 481 -273
rect 501 -275 503 -273
rect 523 -275 525 -273
rect 626 -266 628 -264
rect 571 -275 573 -273
rect 593 -275 595 -273
rect 615 -275 617 -273
<< ntiect1 >>
rect -687 147 -685 149
rect -675 147 -673 149
rect -661 147 -659 149
rect -649 147 -647 149
rect -639 147 -637 149
rect -585 147 -583 149
rect -459 147 -457 149
rect -402 147 -400 149
rect -390 147 -388 149
rect -376 147 -374 149
rect -364 147 -362 149
rect -354 147 -352 149
rect -300 147 -298 149
rect -174 147 -172 149
rect -117 147 -115 149
rect -105 147 -103 149
rect -91 147 -89 149
rect -79 147 -77 149
rect -69 147 -67 149
rect -15 147 -13 149
rect 111 147 113 149
rect 168 147 170 149
rect 180 147 182 149
rect 194 147 196 149
rect 206 147 208 149
rect 216 147 218 149
rect 270 147 272 149
rect 396 147 398 149
rect 501 147 503 149
rect 561 147 563 149
rect 583 147 585 149
rect 595 147 597 149
rect -687 135 -685 137
rect -675 135 -673 137
rect -661 135 -659 137
rect -649 135 -647 137
rect -639 135 -637 137
rect -585 135 -583 137
rect -459 135 -457 137
rect -402 135 -400 137
rect -390 135 -388 137
rect -376 135 -374 137
rect -364 135 -362 137
rect -354 135 -352 137
rect -300 135 -298 137
rect -174 135 -172 137
rect -117 135 -115 137
rect -105 135 -103 137
rect -91 135 -89 137
rect -79 135 -77 137
rect -69 135 -67 137
rect -15 135 -13 137
rect 111 135 113 137
rect 168 135 170 137
rect 180 135 182 137
rect 194 135 196 137
rect 206 135 208 137
rect 216 135 218 137
rect 270 135 272 137
rect 396 135 398 137
rect 501 135 503 137
rect 561 135 563 137
rect 583 135 585 137
rect 595 135 597 137
rect -687 -203 -685 -201
rect -675 -203 -673 -201
rect -661 -203 -659 -201
rect -649 -203 -647 -201
rect -639 -203 -637 -201
rect -585 -203 -583 -201
rect -459 -203 -457 -201
rect -402 -203 -400 -201
rect -390 -203 -388 -201
rect -376 -203 -374 -201
rect -364 -203 -362 -201
rect -354 -203 -352 -201
rect -300 -203 -298 -201
rect -174 -203 -172 -201
rect -117 -203 -115 -201
rect -105 -203 -103 -201
rect -91 -203 -89 -201
rect -79 -203 -77 -201
rect -69 -203 -67 -201
rect -15 -203 -13 -201
rect 111 -203 113 -201
rect 168 -203 170 -201
rect 180 -203 182 -201
rect 194 -203 196 -201
rect 206 -203 208 -201
rect 216 -203 218 -201
rect 270 -203 272 -201
rect 396 -203 398 -201
rect 533 -203 535 -201
rect 625 -203 627 -201
rect -687 -215 -685 -213
rect -675 -215 -673 -213
rect -661 -215 -659 -213
rect -649 -215 -647 -213
rect -639 -215 -637 -213
rect -585 -215 -583 -213
rect -459 -215 -457 -213
rect -402 -215 -400 -213
rect -390 -215 -388 -213
rect -376 -215 -374 -213
rect -364 -215 -362 -213
rect -354 -215 -352 -213
rect -300 -215 -298 -213
rect -174 -215 -172 -213
rect -117 -215 -115 -213
rect -105 -215 -103 -213
rect -91 -215 -89 -213
rect -79 -215 -77 -213
rect -69 -215 -67 -213
rect -15 -215 -13 -213
rect 111 -215 113 -213
rect 168 -215 170 -213
rect 180 -215 182 -213
rect 194 -215 196 -213
rect 206 -215 208 -213
rect 216 -215 218 -213
rect 270 -215 272 -213
rect 396 -215 398 -213
rect 533 -215 535 -213
rect 625 -215 627 -213
<< ptiect1 >>
rect -687 207 -685 209
rect -675 207 -673 209
rect -661 207 -659 209
rect -649 207 -647 209
rect -595 207 -593 209
rect -541 207 -539 209
rect -527 207 -525 209
rect -492 207 -490 209
rect -415 207 -413 209
rect -402 207 -400 209
rect -390 207 -388 209
rect -376 207 -374 209
rect -364 207 -362 209
rect -310 207 -308 209
rect -256 207 -254 209
rect -242 207 -240 209
rect -207 207 -205 209
rect -130 207 -128 209
rect -117 207 -115 209
rect -105 207 -103 209
rect -91 207 -89 209
rect -79 207 -77 209
rect -25 207 -23 209
rect 29 207 31 209
rect 43 207 45 209
rect 78 207 80 209
rect 155 207 157 209
rect 168 207 170 209
rect 180 207 182 209
rect 194 207 196 209
rect 206 207 208 209
rect 260 207 262 209
rect 314 207 316 209
rect 328 207 330 209
rect 363 207 365 209
rect 440 207 442 209
rect 457 207 459 209
rect 517 207 519 209
rect 583 207 585 209
rect 595 207 597 209
rect -687 75 -685 77
rect -675 75 -673 77
rect -661 75 -659 77
rect -649 75 -647 77
rect -595 75 -593 77
rect -541 75 -539 77
rect -527 75 -525 77
rect -492 75 -490 77
rect -415 75 -413 77
rect -402 75 -400 77
rect -390 75 -388 77
rect -376 75 -374 77
rect -364 75 -362 77
rect -310 75 -308 77
rect -256 75 -254 77
rect -242 75 -240 77
rect -207 75 -205 77
rect -130 75 -128 77
rect -117 75 -115 77
rect -105 75 -103 77
rect -91 75 -89 77
rect -79 75 -77 77
rect -25 75 -23 77
rect 29 75 31 77
rect 43 75 45 77
rect 78 75 80 77
rect 155 75 157 77
rect 168 75 170 77
rect 180 75 182 77
rect 194 75 196 77
rect 206 75 208 77
rect 260 75 262 77
rect 314 75 316 77
rect 328 75 330 77
rect 363 75 365 77
rect 440 75 442 77
rect 457 75 459 77
rect 517 75 519 77
rect 583 75 585 77
rect 595 75 597 77
rect -687 -143 -685 -141
rect -675 -143 -673 -141
rect -661 -143 -659 -141
rect -649 -143 -647 -141
rect -595 -143 -593 -141
rect -541 -143 -539 -141
rect -527 -143 -525 -141
rect -492 -143 -490 -141
rect -415 -143 -413 -141
rect -402 -143 -400 -141
rect -390 -143 -388 -141
rect -376 -143 -374 -141
rect -364 -143 -362 -141
rect -310 -143 -308 -141
rect -256 -143 -254 -141
rect -242 -143 -240 -141
rect -207 -143 -205 -141
rect -130 -143 -128 -141
rect -117 -143 -115 -141
rect -105 -143 -103 -141
rect -91 -143 -89 -141
rect -79 -143 -77 -141
rect -25 -143 -23 -141
rect 29 -143 31 -141
rect 43 -143 45 -141
rect 78 -143 80 -141
rect 155 -143 157 -141
rect 168 -143 170 -141
rect 180 -143 182 -141
rect 194 -143 196 -141
rect 206 -143 208 -141
rect 260 -143 262 -141
rect 314 -143 316 -141
rect 328 -143 330 -141
rect 363 -143 365 -141
rect 440 -143 442 -141
rect 461 -143 463 -141
rect 469 -143 471 -141
rect 553 -143 555 -141
rect 561 -143 563 -141
rect -687 -275 -685 -273
rect -675 -275 -673 -273
rect -661 -275 -659 -273
rect -649 -275 -647 -273
rect -595 -275 -593 -273
rect -541 -275 -539 -273
rect -527 -275 -525 -273
rect -492 -275 -490 -273
rect -415 -275 -413 -273
rect -402 -275 -400 -273
rect -390 -275 -388 -273
rect -376 -275 -374 -273
rect -364 -275 -362 -273
rect -310 -275 -308 -273
rect -256 -275 -254 -273
rect -242 -275 -240 -273
rect -207 -275 -205 -273
rect -130 -275 -128 -273
rect -117 -275 -115 -273
rect -105 -275 -103 -273
rect -91 -275 -89 -273
rect -79 -275 -77 -273
rect -25 -275 -23 -273
rect 29 -275 31 -273
rect 43 -275 45 -273
rect 78 -275 80 -273
rect 155 -275 157 -273
rect 168 -275 170 -273
rect 180 -275 182 -273
rect 194 -275 196 -273
rect 206 -275 208 -273
rect 260 -275 262 -273
rect 314 -275 316 -273
rect 328 -275 330 -273
rect 363 -275 365 -273
rect 440 -275 442 -273
rect 461 -275 463 -273
rect 469 -275 471 -273
rect 553 -275 555 -273
rect 561 -275 563 -273
<< pdifct0 >>
rect -685 157 -683 159
rect -659 157 -657 159
rect -636 166 -634 168
rect -636 159 -634 161
rect -614 165 -612 167
rect -614 158 -612 160
rect -604 158 -602 160
rect -582 166 -580 168
rect -582 159 -580 161
rect -560 165 -558 167
rect -560 158 -558 160
rect -550 158 -548 160
rect -528 157 -526 159
rect -528 150 -526 152
rect -493 157 -491 159
rect -493 150 -491 152
rect -456 166 -454 168
rect -456 159 -454 161
rect -434 165 -432 167
rect -434 158 -432 160
rect -424 158 -422 160
rect -400 157 -398 159
rect -374 157 -372 159
rect -351 166 -349 168
rect -351 159 -349 161
rect -329 165 -327 167
rect -329 158 -327 160
rect -319 158 -317 160
rect -297 166 -295 168
rect -297 159 -295 161
rect -275 165 -273 167
rect -275 158 -273 160
rect -265 158 -263 160
rect -243 157 -241 159
rect -243 150 -241 152
rect -208 157 -206 159
rect -208 150 -206 152
rect -171 166 -169 168
rect -171 159 -169 161
rect -149 165 -147 167
rect -149 158 -147 160
rect -139 158 -137 160
rect -115 157 -113 159
rect -89 157 -87 159
rect -66 166 -64 168
rect -66 159 -64 161
rect -44 165 -42 167
rect -44 158 -42 160
rect -34 158 -32 160
rect -12 166 -10 168
rect -12 159 -10 161
rect 10 165 12 167
rect 10 158 12 160
rect 20 158 22 160
rect 42 157 44 159
rect 42 150 44 152
rect 77 157 79 159
rect 77 150 79 152
rect 114 166 116 168
rect 114 159 116 161
rect 136 165 138 167
rect 136 158 138 160
rect 146 158 148 160
rect 170 157 172 159
rect 196 157 198 159
rect 219 166 221 168
rect 219 159 221 161
rect 241 165 243 167
rect 241 158 243 160
rect 251 158 253 160
rect 273 166 275 168
rect 273 159 275 161
rect 295 165 297 167
rect 295 158 297 160
rect 305 158 307 160
rect 327 157 329 159
rect 327 150 329 152
rect 362 157 364 159
rect 362 150 364 152
rect 399 166 401 168
rect 399 159 401 161
rect 421 165 423 167
rect 421 158 423 160
rect 431 158 433 160
rect 466 158 468 160
rect 476 165 478 167
rect 476 158 478 160
rect 498 166 500 168
rect 498 159 500 161
rect 526 158 528 160
rect 536 165 538 167
rect 536 158 538 160
rect 558 166 560 168
rect 558 159 560 161
rect 593 157 595 159
rect -685 125 -683 127
rect -659 125 -657 127
rect -636 123 -634 125
rect -636 116 -634 118
rect -614 124 -612 126
rect -614 117 -612 119
rect -604 124 -602 126
rect -528 132 -526 134
rect -582 123 -580 125
rect -582 116 -580 118
rect -560 124 -558 126
rect -560 117 -558 119
rect -550 124 -548 126
rect -528 125 -526 127
rect -493 132 -491 134
rect -493 125 -491 127
rect -456 123 -454 125
rect -456 116 -454 118
rect -434 124 -432 126
rect -434 117 -432 119
rect -424 124 -422 126
rect -400 125 -398 127
rect -374 125 -372 127
rect -351 123 -349 125
rect -351 116 -349 118
rect -329 124 -327 126
rect -329 117 -327 119
rect -319 124 -317 126
rect -243 132 -241 134
rect -297 123 -295 125
rect -297 116 -295 118
rect -275 124 -273 126
rect -275 117 -273 119
rect -265 124 -263 126
rect -243 125 -241 127
rect -208 132 -206 134
rect -208 125 -206 127
rect -171 123 -169 125
rect -171 116 -169 118
rect -149 124 -147 126
rect -149 117 -147 119
rect -139 124 -137 126
rect -115 125 -113 127
rect -89 125 -87 127
rect -66 123 -64 125
rect -66 116 -64 118
rect -44 124 -42 126
rect -44 117 -42 119
rect -34 124 -32 126
rect 42 132 44 134
rect -12 123 -10 125
rect -12 116 -10 118
rect 10 124 12 126
rect 10 117 12 119
rect 20 124 22 126
rect 42 125 44 127
rect 77 132 79 134
rect 77 125 79 127
rect 114 123 116 125
rect 114 116 116 118
rect 136 124 138 126
rect 136 117 138 119
rect 146 124 148 126
rect 170 125 172 127
rect 196 125 198 127
rect 219 123 221 125
rect 219 116 221 118
rect 241 124 243 126
rect 241 117 243 119
rect 251 124 253 126
rect 327 132 329 134
rect 273 123 275 125
rect 273 116 275 118
rect 295 124 297 126
rect 295 117 297 119
rect 305 124 307 126
rect 327 125 329 127
rect 362 132 364 134
rect 362 125 364 127
rect 399 123 401 125
rect 399 116 401 118
rect 421 124 423 126
rect 421 117 423 119
rect 431 124 433 126
rect 466 124 468 126
rect 476 124 478 126
rect 476 117 478 119
rect 498 123 500 125
rect 498 116 500 118
rect 526 124 528 126
rect 536 124 538 126
rect 536 117 538 119
rect 558 123 560 125
rect 558 116 560 118
rect 593 125 595 127
rect -685 -193 -683 -191
rect -659 -193 -657 -191
rect -636 -184 -634 -182
rect -636 -191 -634 -189
rect -614 -185 -612 -183
rect -614 -192 -612 -190
rect -604 -192 -602 -190
rect -582 -184 -580 -182
rect -582 -191 -580 -189
rect -560 -185 -558 -183
rect -560 -192 -558 -190
rect -550 -192 -548 -190
rect -528 -193 -526 -191
rect -528 -200 -526 -198
rect -493 -193 -491 -191
rect -493 -200 -491 -198
rect -456 -184 -454 -182
rect -456 -191 -454 -189
rect -434 -185 -432 -183
rect -434 -192 -432 -190
rect -424 -192 -422 -190
rect -400 -193 -398 -191
rect -374 -193 -372 -191
rect -351 -184 -349 -182
rect -351 -191 -349 -189
rect -329 -185 -327 -183
rect -329 -192 -327 -190
rect -319 -192 -317 -190
rect -297 -184 -295 -182
rect -297 -191 -295 -189
rect -275 -185 -273 -183
rect -275 -192 -273 -190
rect -265 -192 -263 -190
rect -243 -193 -241 -191
rect -243 -200 -241 -198
rect -208 -193 -206 -191
rect -208 -200 -206 -198
rect -171 -184 -169 -182
rect -171 -191 -169 -189
rect -149 -185 -147 -183
rect -149 -192 -147 -190
rect -139 -192 -137 -190
rect -115 -193 -113 -191
rect -89 -193 -87 -191
rect -66 -184 -64 -182
rect -66 -191 -64 -189
rect -44 -185 -42 -183
rect -44 -192 -42 -190
rect -34 -192 -32 -190
rect -12 -184 -10 -182
rect -12 -191 -10 -189
rect 10 -185 12 -183
rect 10 -192 12 -190
rect 20 -192 22 -190
rect 42 -193 44 -191
rect 42 -200 44 -198
rect 77 -193 79 -191
rect 77 -200 79 -198
rect 114 -184 116 -182
rect 114 -191 116 -189
rect 136 -185 138 -183
rect 136 -192 138 -190
rect 146 -192 148 -190
rect 170 -193 172 -191
rect 196 -193 198 -191
rect 219 -184 221 -182
rect 219 -191 221 -189
rect 241 -185 243 -183
rect 241 -192 243 -190
rect 251 -192 253 -190
rect 273 -184 275 -182
rect 273 -191 275 -189
rect 295 -185 297 -183
rect 295 -192 297 -190
rect 305 -192 307 -190
rect 327 -193 329 -191
rect 327 -200 329 -198
rect 362 -193 364 -191
rect 362 -200 364 -198
rect 399 -184 401 -182
rect 399 -191 401 -189
rect 421 -185 423 -183
rect 421 -192 423 -190
rect 431 -192 433 -190
rect 460 -198 462 -196
rect 491 -193 493 -191
rect 523 -200 525 -198
rect 552 -198 554 -196
rect 583 -193 585 -191
rect 615 -200 617 -198
rect -685 -225 -683 -223
rect -659 -225 -657 -223
rect -636 -227 -634 -225
rect -636 -234 -634 -232
rect -614 -226 -612 -224
rect -614 -233 -612 -231
rect -604 -226 -602 -224
rect -528 -218 -526 -216
rect -582 -227 -580 -225
rect -582 -234 -580 -232
rect -560 -226 -558 -224
rect -560 -233 -558 -231
rect -550 -226 -548 -224
rect -528 -225 -526 -223
rect -493 -218 -491 -216
rect -493 -225 -491 -223
rect -456 -227 -454 -225
rect -456 -234 -454 -232
rect -434 -226 -432 -224
rect -434 -233 -432 -231
rect -424 -226 -422 -224
rect -400 -225 -398 -223
rect -374 -225 -372 -223
rect -351 -227 -349 -225
rect -351 -234 -349 -232
rect -329 -226 -327 -224
rect -329 -233 -327 -231
rect -319 -226 -317 -224
rect -243 -218 -241 -216
rect -297 -227 -295 -225
rect -297 -234 -295 -232
rect -275 -226 -273 -224
rect -275 -233 -273 -231
rect -265 -226 -263 -224
rect -243 -225 -241 -223
rect -208 -218 -206 -216
rect -208 -225 -206 -223
rect -171 -227 -169 -225
rect -171 -234 -169 -232
rect -149 -226 -147 -224
rect -149 -233 -147 -231
rect -139 -226 -137 -224
rect -115 -225 -113 -223
rect -89 -225 -87 -223
rect -66 -227 -64 -225
rect -66 -234 -64 -232
rect -44 -226 -42 -224
rect -44 -233 -42 -231
rect -34 -226 -32 -224
rect 42 -218 44 -216
rect -12 -227 -10 -225
rect -12 -234 -10 -232
rect 10 -226 12 -224
rect 10 -233 12 -231
rect 20 -226 22 -224
rect 42 -225 44 -223
rect 77 -218 79 -216
rect 77 -225 79 -223
rect 114 -227 116 -225
rect 114 -234 116 -232
rect 136 -226 138 -224
rect 136 -233 138 -231
rect 146 -226 148 -224
rect 170 -225 172 -223
rect 196 -225 198 -223
rect 219 -227 221 -225
rect 219 -234 221 -232
rect 241 -226 243 -224
rect 241 -233 243 -231
rect 251 -226 253 -224
rect 327 -218 329 -216
rect 273 -227 275 -225
rect 273 -234 275 -232
rect 295 -226 297 -224
rect 295 -233 297 -231
rect 305 -226 307 -224
rect 327 -225 329 -223
rect 362 -218 364 -216
rect 362 -225 364 -223
rect 460 -220 462 -218
rect 399 -227 401 -225
rect 399 -234 401 -232
rect 421 -226 423 -224
rect 421 -233 423 -231
rect 431 -226 433 -224
rect 491 -225 493 -223
rect 523 -218 525 -216
rect 552 -220 554 -218
rect 583 -225 585 -223
rect 615 -218 617 -216
<< pdifct1 >>
rect -674 172 -672 174
rect -674 165 -672 167
rect -648 172 -646 174
rect -648 165 -646 167
rect -594 170 -592 172
rect -594 163 -592 165
rect -540 170 -538 172
rect -540 163 -538 165
rect -625 147 -623 149
rect -571 147 -569 149
rect -509 164 -507 166
rect -509 157 -507 159
rect -474 164 -472 166
rect -474 157 -472 159
rect -414 170 -412 172
rect -414 163 -412 165
rect -389 172 -387 174
rect -389 165 -387 167
rect -363 172 -361 174
rect -363 165 -361 167
rect -309 170 -307 172
rect -309 163 -307 165
rect -445 147 -443 149
rect -255 170 -253 172
rect -255 163 -253 165
rect -340 147 -338 149
rect -286 147 -284 149
rect -224 164 -222 166
rect -224 157 -222 159
rect -189 164 -187 166
rect -189 157 -187 159
rect -129 170 -127 172
rect -129 163 -127 165
rect -104 172 -102 174
rect -104 165 -102 167
rect -78 172 -76 174
rect -78 165 -76 167
rect -24 170 -22 172
rect -24 163 -22 165
rect -160 147 -158 149
rect 30 170 32 172
rect 30 163 32 165
rect -55 147 -53 149
rect -1 147 1 149
rect 61 164 63 166
rect 61 157 63 159
rect 96 164 98 166
rect 96 157 98 159
rect 156 170 158 172
rect 156 163 158 165
rect 181 172 183 174
rect 181 165 183 167
rect 207 172 209 174
rect 207 165 209 167
rect 261 170 263 172
rect 261 163 263 165
rect 125 147 127 149
rect 315 170 317 172
rect 315 163 317 165
rect 230 147 232 149
rect 284 147 286 149
rect 346 164 348 166
rect 346 157 348 159
rect 381 164 383 166
rect 381 157 383 159
rect 441 170 443 172
rect 441 163 443 165
rect 456 170 458 172
rect 456 163 458 165
rect 516 170 518 172
rect 516 163 518 165
rect 410 147 412 149
rect 582 172 584 174
rect 582 165 584 167
rect 487 147 489 149
rect 547 147 549 149
rect -625 135 -623 137
rect -571 135 -569 137
rect -674 117 -672 119
rect -674 110 -672 112
rect -648 117 -646 119
rect -648 110 -646 112
rect -594 119 -592 121
rect -594 112 -592 114
rect -540 119 -538 121
rect -540 112 -538 114
rect -509 125 -507 127
rect -509 118 -507 120
rect -445 135 -443 137
rect -340 135 -338 137
rect -474 125 -472 127
rect -474 118 -472 120
rect -414 119 -412 121
rect -414 112 -412 114
rect -286 135 -284 137
rect -389 117 -387 119
rect -389 110 -387 112
rect -363 117 -361 119
rect -363 110 -361 112
rect -309 119 -307 121
rect -309 112 -307 114
rect -255 119 -253 121
rect -255 112 -253 114
rect -224 125 -222 127
rect -224 118 -222 120
rect -160 135 -158 137
rect -55 135 -53 137
rect -189 125 -187 127
rect -189 118 -187 120
rect -129 119 -127 121
rect -129 112 -127 114
rect -1 135 1 137
rect -104 117 -102 119
rect -104 110 -102 112
rect -78 117 -76 119
rect -78 110 -76 112
rect -24 119 -22 121
rect -24 112 -22 114
rect 30 119 32 121
rect 30 112 32 114
rect 61 125 63 127
rect 61 118 63 120
rect 125 135 127 137
rect 230 135 232 137
rect 96 125 98 127
rect 96 118 98 120
rect 156 119 158 121
rect 156 112 158 114
rect 284 135 286 137
rect 181 117 183 119
rect 181 110 183 112
rect 207 117 209 119
rect 207 110 209 112
rect 261 119 263 121
rect 261 112 263 114
rect 315 119 317 121
rect 315 112 317 114
rect 346 125 348 127
rect 346 118 348 120
rect 410 135 412 137
rect 487 135 489 137
rect 547 135 549 137
rect 381 125 383 127
rect 381 118 383 120
rect 441 119 443 121
rect 441 112 443 114
rect 456 119 458 121
rect 456 112 458 114
rect 516 119 518 121
rect 516 112 518 114
rect 582 117 584 119
rect 582 110 584 112
rect -674 -178 -672 -176
rect -674 -185 -672 -183
rect -648 -178 -646 -176
rect -648 -185 -646 -183
rect -594 -180 -592 -178
rect -594 -187 -592 -185
rect -540 -180 -538 -178
rect -540 -187 -538 -185
rect -625 -203 -623 -201
rect -571 -203 -569 -201
rect -509 -186 -507 -184
rect -509 -193 -507 -191
rect -474 -186 -472 -184
rect -474 -193 -472 -191
rect -414 -180 -412 -178
rect -414 -187 -412 -185
rect -389 -178 -387 -176
rect -389 -185 -387 -183
rect -363 -178 -361 -176
rect -363 -185 -361 -183
rect -309 -180 -307 -178
rect -309 -187 -307 -185
rect -445 -203 -443 -201
rect -255 -180 -253 -178
rect -255 -187 -253 -185
rect -340 -203 -338 -201
rect -286 -203 -284 -201
rect -224 -186 -222 -184
rect -224 -193 -222 -191
rect -189 -186 -187 -184
rect -189 -193 -187 -191
rect -129 -180 -127 -178
rect -129 -187 -127 -185
rect -104 -178 -102 -176
rect -104 -185 -102 -183
rect -78 -178 -76 -176
rect -78 -185 -76 -183
rect -24 -180 -22 -178
rect -24 -187 -22 -185
rect -160 -203 -158 -201
rect 30 -180 32 -178
rect 30 -187 32 -185
rect -55 -203 -53 -201
rect -1 -203 1 -201
rect 61 -186 63 -184
rect 61 -193 63 -191
rect 96 -186 98 -184
rect 96 -193 98 -191
rect 156 -180 158 -178
rect 156 -187 158 -185
rect 181 -178 183 -176
rect 181 -185 183 -183
rect 207 -178 209 -176
rect 207 -185 209 -183
rect 261 -180 263 -178
rect 261 -187 263 -185
rect 125 -203 127 -201
rect 315 -180 317 -178
rect 315 -187 317 -185
rect 230 -203 232 -201
rect 284 -203 286 -201
rect 346 -186 348 -184
rect 346 -193 348 -191
rect 381 -186 383 -184
rect 381 -193 383 -191
rect 441 -180 443 -178
rect 441 -187 443 -185
rect 534 -178 536 -176
rect 534 -185 536 -183
rect 410 -203 412 -201
rect 626 -178 628 -176
rect 626 -185 628 -183
rect -625 -215 -623 -213
rect -571 -215 -569 -213
rect -674 -233 -672 -231
rect -674 -240 -672 -238
rect -648 -233 -646 -231
rect -648 -240 -646 -238
rect -594 -231 -592 -229
rect -594 -238 -592 -236
rect -540 -231 -538 -229
rect -540 -238 -538 -236
rect -509 -225 -507 -223
rect -509 -232 -507 -230
rect -445 -215 -443 -213
rect -340 -215 -338 -213
rect -474 -225 -472 -223
rect -474 -232 -472 -230
rect -414 -231 -412 -229
rect -414 -238 -412 -236
rect -286 -215 -284 -213
rect -389 -233 -387 -231
rect -389 -240 -387 -238
rect -363 -233 -361 -231
rect -363 -240 -361 -238
rect -309 -231 -307 -229
rect -309 -238 -307 -236
rect -255 -231 -253 -229
rect -255 -238 -253 -236
rect -224 -225 -222 -223
rect -224 -232 -222 -230
rect -160 -215 -158 -213
rect -55 -215 -53 -213
rect -189 -225 -187 -223
rect -189 -232 -187 -230
rect -129 -231 -127 -229
rect -129 -238 -127 -236
rect -1 -215 1 -213
rect -104 -233 -102 -231
rect -104 -240 -102 -238
rect -78 -233 -76 -231
rect -78 -240 -76 -238
rect -24 -231 -22 -229
rect -24 -238 -22 -236
rect 30 -231 32 -229
rect 30 -238 32 -236
rect 61 -225 63 -223
rect 61 -232 63 -230
rect 125 -215 127 -213
rect 230 -215 232 -213
rect 96 -225 98 -223
rect 96 -232 98 -230
rect 156 -231 158 -229
rect 156 -238 158 -236
rect 284 -215 286 -213
rect 181 -233 183 -231
rect 181 -240 183 -238
rect 207 -233 209 -231
rect 207 -240 209 -238
rect 261 -231 263 -229
rect 261 -238 263 -236
rect 315 -231 317 -229
rect 315 -238 317 -236
rect 346 -225 348 -223
rect 346 -232 348 -230
rect 410 -215 412 -213
rect 381 -225 383 -223
rect 381 -232 383 -230
rect 441 -231 443 -229
rect 441 -238 443 -236
rect 534 -233 536 -231
rect 534 -240 536 -238
rect 626 -233 628 -231
rect 626 -240 628 -238
<< alu0 >>
rect -689 195 -685 206
rect -689 193 -688 195
rect -686 193 -685 195
rect -689 191 -685 193
rect -675 188 -674 194
rect -663 195 -659 206
rect -663 193 -662 195
rect -660 193 -659 195
rect -663 191 -659 193
rect -649 188 -648 194
rect -633 200 -603 201
rect -633 198 -631 200
rect -629 198 -603 200
rect -633 197 -603 198
rect -607 193 -603 197
rect -675 169 -674 176
rect -649 169 -648 176
rect -607 189 -598 193
rect -595 189 -594 195
rect -579 200 -549 201
rect -579 198 -577 200
rect -575 198 -549 200
rect -579 197 -549 198
rect -553 193 -549 197
rect -602 183 -598 189
rect -602 181 -601 183
rect -599 181 -598 183
rect -623 176 -617 177
rect -602 176 -598 181
rect -610 172 -598 176
rect -638 168 -632 169
rect -638 166 -636 168
rect -634 166 -632 168
rect -638 161 -632 166
rect -610 169 -606 172
rect -615 167 -606 169
rect -595 168 -594 174
rect -553 189 -544 193
rect -541 189 -540 195
rect -529 197 -525 206
rect -529 195 -528 197
rect -526 195 -525 197
rect -529 193 -525 195
rect -548 183 -544 189
rect -548 181 -547 183
rect -545 181 -544 183
rect -569 176 -563 177
rect -548 176 -544 181
rect -556 172 -544 176
rect -615 165 -614 167
rect -612 165 -606 167
rect -687 159 -681 160
rect -687 157 -685 159
rect -683 157 -681 159
rect -687 150 -681 157
rect -661 159 -655 160
rect -661 157 -659 159
rect -657 157 -655 159
rect -661 150 -655 157
rect -638 159 -636 161
rect -634 160 -632 161
rect -615 160 -611 165
rect -634 159 -614 160
rect -638 158 -614 159
rect -612 158 -611 160
rect -638 156 -611 158
rect -606 160 -600 161
rect -606 158 -604 160
rect -602 158 -600 160
rect -606 150 -600 158
rect -584 168 -578 169
rect -584 166 -582 168
rect -580 166 -578 168
rect -584 161 -578 166
rect -556 169 -552 172
rect -561 167 -552 169
rect -541 168 -540 174
rect -494 197 -490 206
rect -453 200 -423 201
rect -453 198 -451 200
rect -449 198 -423 200
rect -453 197 -423 198
rect -494 195 -493 197
rect -491 195 -490 197
rect -494 193 -490 195
rect -427 193 -423 197
rect -561 165 -560 167
rect -558 165 -552 167
rect -427 189 -418 193
rect -415 189 -414 195
rect -404 195 -400 206
rect -404 193 -403 195
rect -401 193 -400 195
rect -404 191 -400 193
rect -422 183 -418 189
rect -422 181 -421 183
rect -419 181 -418 183
rect -443 176 -437 177
rect -422 176 -418 181
rect -430 172 -418 176
rect -584 159 -582 161
rect -580 160 -578 161
rect -561 160 -557 165
rect -580 159 -560 160
rect -584 158 -560 159
rect -558 158 -557 160
rect -584 156 -557 158
rect -552 160 -546 161
rect -552 158 -550 160
rect -548 158 -546 160
rect -552 150 -546 158
rect -458 168 -452 169
rect -458 166 -456 168
rect -454 166 -452 168
rect -529 159 -525 161
rect -529 157 -528 159
rect -526 157 -525 159
rect -529 152 -525 157
rect -494 159 -490 161
rect -494 157 -493 159
rect -491 157 -490 159
rect -529 150 -528 152
rect -526 150 -525 152
rect -494 152 -490 157
rect -458 161 -452 166
rect -430 169 -426 172
rect -435 167 -426 169
rect -415 168 -414 174
rect -390 188 -389 194
rect -378 195 -374 206
rect -378 193 -377 195
rect -375 193 -374 195
rect -378 191 -374 193
rect -364 188 -363 194
rect -348 200 -318 201
rect -348 198 -346 200
rect -344 198 -318 200
rect -348 197 -318 198
rect -322 193 -318 197
rect -390 169 -389 176
rect -364 169 -363 176
rect -322 189 -313 193
rect -310 189 -309 195
rect -294 200 -264 201
rect -294 198 -292 200
rect -290 198 -264 200
rect -294 197 -264 198
rect -268 193 -264 197
rect -317 183 -313 189
rect -317 181 -316 183
rect -314 181 -313 183
rect -338 176 -332 177
rect -317 176 -313 181
rect -325 172 -313 176
rect -435 165 -434 167
rect -432 165 -426 167
rect -458 159 -456 161
rect -454 160 -452 161
rect -435 160 -431 165
rect -353 168 -347 169
rect -353 166 -351 168
rect -349 166 -347 168
rect -454 159 -434 160
rect -458 158 -434 159
rect -432 158 -431 160
rect -458 156 -431 158
rect -426 160 -420 161
rect -426 158 -424 160
rect -422 158 -420 160
rect -494 150 -493 152
rect -491 150 -490 152
rect -426 150 -420 158
rect -353 161 -347 166
rect -325 169 -321 172
rect -330 167 -321 169
rect -310 168 -309 174
rect -268 189 -259 193
rect -256 189 -255 195
rect -244 197 -240 206
rect -244 195 -243 197
rect -241 195 -240 197
rect -244 193 -240 195
rect -263 183 -259 189
rect -263 181 -262 183
rect -260 181 -259 183
rect -284 176 -278 177
rect -263 176 -259 181
rect -271 172 -259 176
rect -330 165 -329 167
rect -327 165 -321 167
rect -402 159 -396 160
rect -402 157 -400 159
rect -398 157 -396 159
rect -402 150 -396 157
rect -376 159 -370 160
rect -376 157 -374 159
rect -372 157 -370 159
rect -376 150 -370 157
rect -353 159 -351 161
rect -349 160 -347 161
rect -330 160 -326 165
rect -349 159 -329 160
rect -353 158 -329 159
rect -327 158 -326 160
rect -353 156 -326 158
rect -321 160 -315 161
rect -321 158 -319 160
rect -317 158 -315 160
rect -321 150 -315 158
rect -299 168 -293 169
rect -299 166 -297 168
rect -295 166 -293 168
rect -299 161 -293 166
rect -271 169 -267 172
rect -276 167 -267 169
rect -256 168 -255 174
rect -209 197 -205 206
rect -168 200 -138 201
rect -168 198 -166 200
rect -164 198 -138 200
rect -168 197 -138 198
rect -209 195 -208 197
rect -206 195 -205 197
rect -209 193 -205 195
rect -142 193 -138 197
rect -276 165 -275 167
rect -273 165 -267 167
rect -142 189 -133 193
rect -130 189 -129 195
rect -119 195 -115 206
rect -119 193 -118 195
rect -116 193 -115 195
rect -119 191 -115 193
rect -137 183 -133 189
rect -137 181 -136 183
rect -134 181 -133 183
rect -158 176 -152 177
rect -137 176 -133 181
rect -145 172 -133 176
rect -299 159 -297 161
rect -295 160 -293 161
rect -276 160 -272 165
rect -295 159 -275 160
rect -299 158 -275 159
rect -273 158 -272 160
rect -299 156 -272 158
rect -267 160 -261 161
rect -267 158 -265 160
rect -263 158 -261 160
rect -267 150 -261 158
rect -173 168 -167 169
rect -173 166 -171 168
rect -169 166 -167 168
rect -244 159 -240 161
rect -244 157 -243 159
rect -241 157 -240 159
rect -244 152 -240 157
rect -209 159 -205 161
rect -209 157 -208 159
rect -206 157 -205 159
rect -244 150 -243 152
rect -241 150 -240 152
rect -209 152 -205 157
rect -173 161 -167 166
rect -145 169 -141 172
rect -150 167 -141 169
rect -130 168 -129 174
rect -105 188 -104 194
rect -93 195 -89 206
rect -93 193 -92 195
rect -90 193 -89 195
rect -93 191 -89 193
rect -79 188 -78 194
rect -63 200 -33 201
rect -63 198 -61 200
rect -59 198 -33 200
rect -63 197 -33 198
rect -37 193 -33 197
rect -105 169 -104 176
rect -79 169 -78 176
rect -37 189 -28 193
rect -25 189 -24 195
rect -9 200 21 201
rect -9 198 -7 200
rect -5 198 21 200
rect -9 197 21 198
rect 17 193 21 197
rect -32 183 -28 189
rect -32 181 -31 183
rect -29 181 -28 183
rect -53 176 -47 177
rect -32 176 -28 181
rect -40 172 -28 176
rect -150 165 -149 167
rect -147 165 -141 167
rect -173 159 -171 161
rect -169 160 -167 161
rect -150 160 -146 165
rect -68 168 -62 169
rect -68 166 -66 168
rect -64 166 -62 168
rect -169 159 -149 160
rect -173 158 -149 159
rect -147 158 -146 160
rect -173 156 -146 158
rect -141 160 -135 161
rect -141 158 -139 160
rect -137 158 -135 160
rect -209 150 -208 152
rect -206 150 -205 152
rect -141 150 -135 158
rect -68 161 -62 166
rect -40 169 -36 172
rect -45 167 -36 169
rect -25 168 -24 174
rect 17 189 26 193
rect 29 189 30 195
rect 41 197 45 206
rect 41 195 42 197
rect 44 195 45 197
rect 41 193 45 195
rect 22 183 26 189
rect 22 181 23 183
rect 25 181 26 183
rect 1 176 7 177
rect 22 176 26 181
rect 14 172 26 176
rect -45 165 -44 167
rect -42 165 -36 167
rect -117 159 -111 160
rect -117 157 -115 159
rect -113 157 -111 159
rect -117 150 -111 157
rect -91 159 -85 160
rect -91 157 -89 159
rect -87 157 -85 159
rect -91 150 -85 157
rect -68 159 -66 161
rect -64 160 -62 161
rect -45 160 -41 165
rect -64 159 -44 160
rect -68 158 -44 159
rect -42 158 -41 160
rect -68 156 -41 158
rect -36 160 -30 161
rect -36 158 -34 160
rect -32 158 -30 160
rect -36 150 -30 158
rect -14 168 -8 169
rect -14 166 -12 168
rect -10 166 -8 168
rect -14 161 -8 166
rect 14 169 18 172
rect 9 167 18 169
rect 29 168 30 174
rect 76 197 80 206
rect 117 200 147 201
rect 117 198 119 200
rect 121 198 147 200
rect 117 197 147 198
rect 76 195 77 197
rect 79 195 80 197
rect 76 193 80 195
rect 143 193 147 197
rect 9 165 10 167
rect 12 165 18 167
rect 143 189 152 193
rect 155 189 156 195
rect 166 195 170 206
rect 166 193 167 195
rect 169 193 170 195
rect 166 191 170 193
rect 148 183 152 189
rect 148 181 149 183
rect 151 181 152 183
rect 127 176 133 177
rect 148 176 152 181
rect 140 172 152 176
rect -14 159 -12 161
rect -10 160 -8 161
rect 9 160 13 165
rect -10 159 10 160
rect -14 158 10 159
rect 12 158 13 160
rect -14 156 13 158
rect 18 160 24 161
rect 18 158 20 160
rect 22 158 24 160
rect 18 150 24 158
rect 112 168 118 169
rect 112 166 114 168
rect 116 166 118 168
rect 41 159 45 161
rect 41 157 42 159
rect 44 157 45 159
rect 41 152 45 157
rect 76 159 80 161
rect 76 157 77 159
rect 79 157 80 159
rect 41 150 42 152
rect 44 150 45 152
rect 76 152 80 157
rect 112 161 118 166
rect 140 169 144 172
rect 135 167 144 169
rect 155 168 156 174
rect 180 188 181 194
rect 192 195 196 206
rect 192 193 193 195
rect 195 193 196 195
rect 192 191 196 193
rect 206 188 207 194
rect 222 200 252 201
rect 222 198 224 200
rect 226 198 252 200
rect 222 197 252 198
rect 248 193 252 197
rect 180 169 181 176
rect 206 169 207 176
rect 248 189 257 193
rect 260 189 261 195
rect 276 200 306 201
rect 276 198 278 200
rect 280 198 306 200
rect 276 197 306 198
rect 302 193 306 197
rect 253 183 257 189
rect 253 181 254 183
rect 256 181 257 183
rect 232 176 238 177
rect 253 176 257 181
rect 245 172 257 176
rect 135 165 136 167
rect 138 165 144 167
rect 112 159 114 161
rect 116 160 118 161
rect 135 160 139 165
rect 217 168 223 169
rect 217 166 219 168
rect 221 166 223 168
rect 116 159 136 160
rect 112 158 136 159
rect 138 158 139 160
rect 112 156 139 158
rect 144 160 150 161
rect 144 158 146 160
rect 148 158 150 160
rect 76 150 77 152
rect 79 150 80 152
rect 144 150 150 158
rect 217 161 223 166
rect 245 169 249 172
rect 240 167 249 169
rect 260 168 261 174
rect 302 189 311 193
rect 314 189 315 195
rect 326 197 330 206
rect 326 195 327 197
rect 329 195 330 197
rect 326 193 330 195
rect 307 183 311 189
rect 307 181 308 183
rect 310 181 311 183
rect 286 176 292 177
rect 307 176 311 181
rect 299 172 311 176
rect 240 165 241 167
rect 243 165 249 167
rect 168 159 174 160
rect 168 157 170 159
rect 172 157 174 159
rect 168 150 174 157
rect 194 159 200 160
rect 194 157 196 159
rect 198 157 200 159
rect 194 150 200 157
rect 217 159 219 161
rect 221 160 223 161
rect 240 160 244 165
rect 221 159 241 160
rect 217 158 241 159
rect 243 158 244 160
rect 217 156 244 158
rect 249 160 255 161
rect 249 158 251 160
rect 253 158 255 160
rect 249 150 255 158
rect 271 168 277 169
rect 271 166 273 168
rect 275 166 277 168
rect 271 161 277 166
rect 299 169 303 172
rect 294 167 303 169
rect 314 168 315 174
rect 361 197 365 206
rect 402 200 432 201
rect 402 198 404 200
rect 406 198 432 200
rect 402 197 432 198
rect 361 195 362 197
rect 364 195 365 197
rect 361 193 365 195
rect 428 193 432 197
rect 294 165 295 167
rect 297 165 303 167
rect 428 189 437 193
rect 440 189 441 195
rect 433 183 437 189
rect 433 181 434 183
rect 436 181 437 183
rect 412 176 418 177
rect 433 176 437 181
rect 425 172 437 176
rect 271 159 273 161
rect 275 160 277 161
rect 294 160 298 165
rect 275 159 295 160
rect 271 158 295 159
rect 297 158 298 160
rect 271 156 298 158
rect 303 160 309 161
rect 303 158 305 160
rect 307 158 309 160
rect 303 150 309 158
rect 397 168 403 169
rect 397 166 399 168
rect 401 166 403 168
rect 326 159 330 161
rect 326 157 327 159
rect 329 157 330 159
rect 326 152 330 157
rect 361 159 365 161
rect 361 157 362 159
rect 364 157 365 159
rect 326 150 327 152
rect 329 150 330 152
rect 361 152 365 157
rect 397 161 403 166
rect 425 169 429 172
rect 420 167 429 169
rect 440 168 441 174
rect 420 165 421 167
rect 423 165 429 167
rect 397 159 399 161
rect 401 160 403 161
rect 420 160 424 165
rect 401 159 421 160
rect 397 158 421 159
rect 423 158 424 160
rect 397 156 424 158
rect 429 160 435 161
rect 429 158 431 160
rect 433 158 435 160
rect 361 150 362 152
rect 364 150 365 152
rect 429 150 435 158
rect 467 200 497 201
rect 467 198 493 200
rect 495 198 497 200
rect 467 197 497 198
rect 458 189 459 195
rect 467 193 471 197
rect 527 200 557 201
rect 527 198 553 200
rect 555 198 557 200
rect 527 197 557 198
rect 462 189 471 193
rect 462 183 466 189
rect 518 189 519 195
rect 527 193 531 197
rect 522 189 531 193
rect 462 181 463 183
rect 465 181 466 183
rect 462 176 466 181
rect 481 176 487 177
rect 458 168 459 174
rect 462 172 474 176
rect 522 183 526 189
rect 522 181 523 183
rect 525 181 526 183
rect 522 176 526 181
rect 595 195 599 206
rect 541 176 547 177
rect 470 169 474 172
rect 470 167 479 169
rect 470 165 476 167
rect 478 165 479 167
rect 464 160 470 161
rect 464 158 466 160
rect 468 158 470 160
rect 464 150 470 158
rect 475 160 479 165
rect 496 168 502 169
rect 496 166 498 168
rect 500 166 502 168
rect 496 161 502 166
rect 496 160 498 161
rect 475 158 476 160
rect 478 159 498 160
rect 500 159 502 161
rect 478 158 502 159
rect 475 156 502 158
rect 518 168 519 174
rect 522 172 534 176
rect 584 188 585 194
rect 595 193 596 195
rect 598 193 599 195
rect 595 191 599 193
rect 530 169 534 172
rect 530 167 539 169
rect 530 165 536 167
rect 538 165 539 167
rect 524 160 530 161
rect 524 158 526 160
rect 528 158 530 160
rect 524 150 530 158
rect 535 160 539 165
rect 584 169 585 176
rect 556 168 562 169
rect 556 166 558 168
rect 560 166 562 168
rect 556 161 562 166
rect 556 160 558 161
rect 535 158 536 160
rect 538 159 558 160
rect 560 159 562 161
rect 538 158 562 159
rect 535 156 562 158
rect 591 159 597 160
rect 591 157 593 159
rect 595 157 597 159
rect 591 150 597 157
rect -687 127 -681 134
rect -687 125 -685 127
rect -683 125 -681 127
rect -687 124 -681 125
rect -661 127 -655 134
rect -661 125 -659 127
rect -657 125 -655 127
rect -661 124 -655 125
rect -638 126 -611 128
rect -638 125 -614 126
rect -638 123 -636 125
rect -634 124 -614 125
rect -612 124 -611 126
rect -634 123 -632 124
rect -638 118 -632 123
rect -638 116 -636 118
rect -634 116 -632 118
rect -638 115 -632 116
rect -675 108 -674 115
rect -689 91 -685 93
rect -649 108 -648 115
rect -615 119 -611 124
rect -606 126 -600 134
rect -606 124 -604 126
rect -602 124 -600 126
rect -606 123 -600 124
rect -615 117 -614 119
rect -612 117 -606 119
rect -615 115 -606 117
rect -610 112 -606 115
rect -689 89 -688 91
rect -686 89 -685 91
rect -675 90 -674 96
rect -689 78 -685 89
rect -663 91 -659 93
rect -610 108 -598 112
rect -595 110 -594 116
rect -584 126 -557 128
rect -584 125 -560 126
rect -584 123 -582 125
rect -580 124 -560 125
rect -558 124 -557 126
rect -580 123 -578 124
rect -584 118 -578 123
rect -584 116 -582 118
rect -580 116 -578 118
rect -584 115 -578 116
rect -561 119 -557 124
rect -552 126 -546 134
rect -529 132 -528 134
rect -526 132 -525 134
rect -552 124 -550 126
rect -548 124 -546 126
rect -552 123 -546 124
rect -529 127 -525 132
rect -494 132 -493 134
rect -491 132 -490 134
rect -529 125 -528 127
rect -526 125 -525 127
rect -529 123 -525 125
rect -561 117 -560 119
rect -558 117 -552 119
rect -561 115 -552 117
rect -494 127 -490 132
rect -494 125 -493 127
rect -491 125 -490 127
rect -494 123 -490 125
rect -458 126 -431 128
rect -458 125 -434 126
rect -458 123 -456 125
rect -454 124 -434 125
rect -432 124 -431 126
rect -454 123 -452 124
rect -556 112 -552 115
rect -623 107 -617 108
rect -663 89 -662 91
rect -660 89 -659 91
rect -649 90 -648 96
rect -663 78 -659 89
rect -602 103 -598 108
rect -602 101 -601 103
rect -599 101 -598 103
rect -602 95 -598 101
rect -556 108 -544 112
rect -541 110 -540 116
rect -569 107 -563 108
rect -607 91 -598 95
rect -607 87 -603 91
rect -595 89 -594 95
rect -548 103 -544 108
rect -548 101 -547 103
rect -545 101 -544 103
rect -548 95 -544 101
rect -553 91 -544 95
rect -633 86 -603 87
rect -633 84 -631 86
rect -629 84 -603 86
rect -633 83 -603 84
rect -553 87 -549 91
rect -541 89 -540 95
rect -579 86 -549 87
rect -579 84 -577 86
rect -575 84 -549 86
rect -579 83 -549 84
rect -529 89 -525 91
rect -458 118 -452 123
rect -458 116 -456 118
rect -454 116 -452 118
rect -458 115 -452 116
rect -435 119 -431 124
rect -426 126 -420 134
rect -426 124 -424 126
rect -422 124 -420 126
rect -426 123 -420 124
rect -402 127 -396 134
rect -402 125 -400 127
rect -398 125 -396 127
rect -402 124 -396 125
rect -376 127 -370 134
rect -376 125 -374 127
rect -372 125 -370 127
rect -376 124 -370 125
rect -353 126 -326 128
rect -353 125 -329 126
rect -353 123 -351 125
rect -349 124 -329 125
rect -327 124 -326 126
rect -349 123 -347 124
rect -435 117 -434 119
rect -432 117 -426 119
rect -435 115 -426 117
rect -430 112 -426 115
rect -430 108 -418 112
rect -415 110 -414 116
rect -353 118 -347 123
rect -353 116 -351 118
rect -349 116 -347 118
rect -353 115 -347 116
rect -443 107 -437 108
rect -422 103 -418 108
rect -422 101 -421 103
rect -419 101 -418 103
rect -422 95 -418 101
rect -390 108 -389 115
rect -427 91 -418 95
rect -529 87 -528 89
rect -526 87 -525 89
rect -529 78 -525 87
rect -494 89 -490 91
rect -494 87 -493 89
rect -491 87 -490 89
rect -427 87 -423 91
rect -415 89 -414 95
rect -494 78 -490 87
rect -453 86 -423 87
rect -453 84 -451 86
rect -449 84 -423 86
rect -453 83 -423 84
rect -404 91 -400 93
rect -364 108 -363 115
rect -330 119 -326 124
rect -321 126 -315 134
rect -321 124 -319 126
rect -317 124 -315 126
rect -321 123 -315 124
rect -330 117 -329 119
rect -327 117 -321 119
rect -330 115 -321 117
rect -325 112 -321 115
rect -404 89 -403 91
rect -401 89 -400 91
rect -390 90 -389 96
rect -404 78 -400 89
rect -378 91 -374 93
rect -325 108 -313 112
rect -310 110 -309 116
rect -299 126 -272 128
rect -299 125 -275 126
rect -299 123 -297 125
rect -295 124 -275 125
rect -273 124 -272 126
rect -295 123 -293 124
rect -299 118 -293 123
rect -299 116 -297 118
rect -295 116 -293 118
rect -299 115 -293 116
rect -276 119 -272 124
rect -267 126 -261 134
rect -244 132 -243 134
rect -241 132 -240 134
rect -267 124 -265 126
rect -263 124 -261 126
rect -267 123 -261 124
rect -244 127 -240 132
rect -209 132 -208 134
rect -206 132 -205 134
rect -244 125 -243 127
rect -241 125 -240 127
rect -244 123 -240 125
rect -276 117 -275 119
rect -273 117 -267 119
rect -276 115 -267 117
rect -209 127 -205 132
rect -209 125 -208 127
rect -206 125 -205 127
rect -209 123 -205 125
rect -173 126 -146 128
rect -173 125 -149 126
rect -173 123 -171 125
rect -169 124 -149 125
rect -147 124 -146 126
rect -169 123 -167 124
rect -271 112 -267 115
rect -338 107 -332 108
rect -378 89 -377 91
rect -375 89 -374 91
rect -364 90 -363 96
rect -378 78 -374 89
rect -317 103 -313 108
rect -317 101 -316 103
rect -314 101 -313 103
rect -317 95 -313 101
rect -271 108 -259 112
rect -256 110 -255 116
rect -284 107 -278 108
rect -322 91 -313 95
rect -322 87 -318 91
rect -310 89 -309 95
rect -263 103 -259 108
rect -263 101 -262 103
rect -260 101 -259 103
rect -263 95 -259 101
rect -268 91 -259 95
rect -348 86 -318 87
rect -348 84 -346 86
rect -344 84 -318 86
rect -348 83 -318 84
rect -268 87 -264 91
rect -256 89 -255 95
rect -294 86 -264 87
rect -294 84 -292 86
rect -290 84 -264 86
rect -294 83 -264 84
rect -244 89 -240 91
rect -173 118 -167 123
rect -173 116 -171 118
rect -169 116 -167 118
rect -173 115 -167 116
rect -150 119 -146 124
rect -141 126 -135 134
rect -141 124 -139 126
rect -137 124 -135 126
rect -141 123 -135 124
rect -117 127 -111 134
rect -117 125 -115 127
rect -113 125 -111 127
rect -117 124 -111 125
rect -91 127 -85 134
rect -91 125 -89 127
rect -87 125 -85 127
rect -91 124 -85 125
rect -68 126 -41 128
rect -68 125 -44 126
rect -68 123 -66 125
rect -64 124 -44 125
rect -42 124 -41 126
rect -64 123 -62 124
rect -150 117 -149 119
rect -147 117 -141 119
rect -150 115 -141 117
rect -145 112 -141 115
rect -145 108 -133 112
rect -130 110 -129 116
rect -68 118 -62 123
rect -68 116 -66 118
rect -64 116 -62 118
rect -68 115 -62 116
rect -158 107 -152 108
rect -137 103 -133 108
rect -137 101 -136 103
rect -134 101 -133 103
rect -137 95 -133 101
rect -105 108 -104 115
rect -142 91 -133 95
rect -244 87 -243 89
rect -241 87 -240 89
rect -244 78 -240 87
rect -209 89 -205 91
rect -209 87 -208 89
rect -206 87 -205 89
rect -142 87 -138 91
rect -130 89 -129 95
rect -209 78 -205 87
rect -168 86 -138 87
rect -168 84 -166 86
rect -164 84 -138 86
rect -168 83 -138 84
rect -119 91 -115 93
rect -79 108 -78 115
rect -45 119 -41 124
rect -36 126 -30 134
rect -36 124 -34 126
rect -32 124 -30 126
rect -36 123 -30 124
rect -45 117 -44 119
rect -42 117 -36 119
rect -45 115 -36 117
rect -40 112 -36 115
rect -119 89 -118 91
rect -116 89 -115 91
rect -105 90 -104 96
rect -119 78 -115 89
rect -93 91 -89 93
rect -40 108 -28 112
rect -25 110 -24 116
rect -14 126 13 128
rect -14 125 10 126
rect -14 123 -12 125
rect -10 124 10 125
rect 12 124 13 126
rect -10 123 -8 124
rect -14 118 -8 123
rect -14 116 -12 118
rect -10 116 -8 118
rect -14 115 -8 116
rect 9 119 13 124
rect 18 126 24 134
rect 41 132 42 134
rect 44 132 45 134
rect 18 124 20 126
rect 22 124 24 126
rect 18 123 24 124
rect 41 127 45 132
rect 76 132 77 134
rect 79 132 80 134
rect 41 125 42 127
rect 44 125 45 127
rect 41 123 45 125
rect 9 117 10 119
rect 12 117 18 119
rect 9 115 18 117
rect 76 127 80 132
rect 76 125 77 127
rect 79 125 80 127
rect 76 123 80 125
rect 112 126 139 128
rect 112 125 136 126
rect 112 123 114 125
rect 116 124 136 125
rect 138 124 139 126
rect 116 123 118 124
rect 14 112 18 115
rect -53 107 -47 108
rect -93 89 -92 91
rect -90 89 -89 91
rect -79 90 -78 96
rect -93 78 -89 89
rect -32 103 -28 108
rect -32 101 -31 103
rect -29 101 -28 103
rect -32 95 -28 101
rect 14 108 26 112
rect 29 110 30 116
rect 1 107 7 108
rect -37 91 -28 95
rect -37 87 -33 91
rect -25 89 -24 95
rect 22 103 26 108
rect 22 101 23 103
rect 25 101 26 103
rect 22 95 26 101
rect 17 91 26 95
rect -63 86 -33 87
rect -63 84 -61 86
rect -59 84 -33 86
rect -63 83 -33 84
rect 17 87 21 91
rect 29 89 30 95
rect -9 86 21 87
rect -9 84 -7 86
rect -5 84 21 86
rect -9 83 21 84
rect 41 89 45 91
rect 112 118 118 123
rect 112 116 114 118
rect 116 116 118 118
rect 112 115 118 116
rect 135 119 139 124
rect 144 126 150 134
rect 144 124 146 126
rect 148 124 150 126
rect 144 123 150 124
rect 168 127 174 134
rect 168 125 170 127
rect 172 125 174 127
rect 168 124 174 125
rect 194 127 200 134
rect 194 125 196 127
rect 198 125 200 127
rect 194 124 200 125
rect 217 126 244 128
rect 217 125 241 126
rect 217 123 219 125
rect 221 124 241 125
rect 243 124 244 126
rect 221 123 223 124
rect 135 117 136 119
rect 138 117 144 119
rect 135 115 144 117
rect 140 112 144 115
rect 140 108 152 112
rect 155 110 156 116
rect 217 118 223 123
rect 217 116 219 118
rect 221 116 223 118
rect 217 115 223 116
rect 127 107 133 108
rect 148 103 152 108
rect 148 101 149 103
rect 151 101 152 103
rect 148 95 152 101
rect 180 108 181 115
rect 143 91 152 95
rect 41 87 42 89
rect 44 87 45 89
rect 41 78 45 87
rect 76 89 80 91
rect 76 87 77 89
rect 79 87 80 89
rect 143 87 147 91
rect 155 89 156 95
rect 76 78 80 87
rect 117 86 147 87
rect 117 84 119 86
rect 121 84 147 86
rect 117 83 147 84
rect 166 91 170 93
rect 206 108 207 115
rect 240 119 244 124
rect 249 126 255 134
rect 249 124 251 126
rect 253 124 255 126
rect 249 123 255 124
rect 240 117 241 119
rect 243 117 249 119
rect 240 115 249 117
rect 245 112 249 115
rect 166 89 167 91
rect 169 89 170 91
rect 180 90 181 96
rect 166 78 170 89
rect 192 91 196 93
rect 245 108 257 112
rect 260 110 261 116
rect 271 126 298 128
rect 271 125 295 126
rect 271 123 273 125
rect 275 124 295 125
rect 297 124 298 126
rect 275 123 277 124
rect 271 118 277 123
rect 271 116 273 118
rect 275 116 277 118
rect 271 115 277 116
rect 294 119 298 124
rect 303 126 309 134
rect 326 132 327 134
rect 329 132 330 134
rect 303 124 305 126
rect 307 124 309 126
rect 303 123 309 124
rect 326 127 330 132
rect 361 132 362 134
rect 364 132 365 134
rect 326 125 327 127
rect 329 125 330 127
rect 326 123 330 125
rect 294 117 295 119
rect 297 117 303 119
rect 294 115 303 117
rect 361 127 365 132
rect 361 125 362 127
rect 364 125 365 127
rect 361 123 365 125
rect 397 126 424 128
rect 397 125 421 126
rect 397 123 399 125
rect 401 124 421 125
rect 423 124 424 126
rect 401 123 403 124
rect 299 112 303 115
rect 232 107 238 108
rect 192 89 193 91
rect 195 89 196 91
rect 206 90 207 96
rect 192 78 196 89
rect 253 103 257 108
rect 253 101 254 103
rect 256 101 257 103
rect 253 95 257 101
rect 299 108 311 112
rect 314 110 315 116
rect 286 107 292 108
rect 248 91 257 95
rect 248 87 252 91
rect 260 89 261 95
rect 307 103 311 108
rect 307 101 308 103
rect 310 101 311 103
rect 307 95 311 101
rect 302 91 311 95
rect 222 86 252 87
rect 222 84 224 86
rect 226 84 252 86
rect 222 83 252 84
rect 302 87 306 91
rect 314 89 315 95
rect 276 86 306 87
rect 276 84 278 86
rect 280 84 306 86
rect 276 83 306 84
rect 326 89 330 91
rect 397 118 403 123
rect 397 116 399 118
rect 401 116 403 118
rect 397 115 403 116
rect 420 119 424 124
rect 429 126 435 134
rect 429 124 431 126
rect 433 124 435 126
rect 429 123 435 124
rect 420 117 421 119
rect 423 117 429 119
rect 420 115 429 117
rect 425 112 429 115
rect 425 108 437 112
rect 440 110 441 116
rect 412 107 418 108
rect 433 103 437 108
rect 433 101 434 103
rect 436 101 437 103
rect 433 95 437 101
rect 428 91 437 95
rect 326 87 327 89
rect 329 87 330 89
rect 326 78 330 87
rect 361 89 365 91
rect 361 87 362 89
rect 364 87 365 89
rect 428 87 432 91
rect 440 89 441 95
rect 361 78 365 87
rect 402 86 432 87
rect 402 84 404 86
rect 406 84 432 86
rect 402 83 432 84
rect 464 126 470 134
rect 464 124 466 126
rect 468 124 470 126
rect 464 123 470 124
rect 475 126 502 128
rect 475 124 476 126
rect 478 125 502 126
rect 478 124 498 125
rect 475 119 479 124
rect 496 123 498 124
rect 500 123 502 125
rect 470 117 476 119
rect 478 117 479 119
rect 458 110 459 116
rect 470 115 479 117
rect 470 112 474 115
rect 496 118 502 123
rect 496 116 498 118
rect 500 116 502 118
rect 496 115 502 116
rect 524 126 530 134
rect 524 124 526 126
rect 528 124 530 126
rect 524 123 530 124
rect 535 126 562 128
rect 535 124 536 126
rect 538 125 562 126
rect 538 124 558 125
rect 535 119 539 124
rect 556 123 558 124
rect 560 123 562 125
rect 591 127 597 134
rect 591 125 593 127
rect 595 125 597 127
rect 591 124 597 125
rect 530 117 536 119
rect 538 117 539 119
rect 462 108 474 112
rect 462 103 466 108
rect 481 107 487 108
rect 462 101 463 103
rect 465 101 466 103
rect 462 95 466 101
rect 458 89 459 95
rect 462 91 471 95
rect 518 110 519 116
rect 530 115 539 117
rect 530 112 534 115
rect 556 118 562 123
rect 556 116 558 118
rect 560 116 562 118
rect 556 115 562 116
rect 522 108 534 112
rect 522 103 526 108
rect 541 107 547 108
rect 522 101 523 103
rect 525 101 526 103
rect 522 95 526 101
rect 467 87 471 91
rect 467 86 497 87
rect 467 84 493 86
rect 495 84 497 86
rect 467 83 497 84
rect 518 89 519 95
rect 522 91 531 95
rect 584 108 585 115
rect 527 87 531 91
rect 584 90 585 96
rect 595 91 599 93
rect 527 86 557 87
rect 527 84 553 86
rect 555 84 557 86
rect 527 83 557 84
rect 595 89 596 91
rect 598 89 599 91
rect 595 78 599 89
rect -689 -155 -685 -144
rect -689 -157 -688 -155
rect -686 -157 -685 -155
rect -689 -159 -685 -157
rect -675 -162 -674 -156
rect -663 -155 -659 -144
rect -663 -157 -662 -155
rect -660 -157 -659 -155
rect -663 -159 -659 -157
rect -649 -162 -648 -156
rect -633 -150 -603 -149
rect -633 -152 -631 -150
rect -629 -152 -603 -150
rect -633 -153 -603 -152
rect -607 -157 -603 -153
rect -675 -181 -674 -174
rect -649 -181 -648 -174
rect -607 -161 -598 -157
rect -595 -161 -594 -155
rect -579 -150 -549 -149
rect -579 -152 -577 -150
rect -575 -152 -549 -150
rect -579 -153 -549 -152
rect -553 -157 -549 -153
rect -602 -167 -598 -161
rect -602 -169 -601 -167
rect -599 -169 -598 -167
rect -623 -174 -617 -173
rect -602 -174 -598 -169
rect -610 -178 -598 -174
rect -638 -182 -632 -181
rect -638 -184 -636 -182
rect -634 -184 -632 -182
rect -638 -189 -632 -184
rect -610 -181 -606 -178
rect -615 -183 -606 -181
rect -595 -182 -594 -176
rect -553 -161 -544 -157
rect -541 -161 -540 -155
rect -529 -153 -525 -144
rect -529 -155 -528 -153
rect -526 -155 -525 -153
rect -529 -157 -525 -155
rect -548 -167 -544 -161
rect -548 -169 -547 -167
rect -545 -169 -544 -167
rect -569 -174 -563 -173
rect -548 -174 -544 -169
rect -556 -178 -544 -174
rect -615 -185 -614 -183
rect -612 -185 -606 -183
rect -687 -191 -681 -190
rect -687 -193 -685 -191
rect -683 -193 -681 -191
rect -687 -200 -681 -193
rect -661 -191 -655 -190
rect -661 -193 -659 -191
rect -657 -193 -655 -191
rect -661 -200 -655 -193
rect -638 -191 -636 -189
rect -634 -190 -632 -189
rect -615 -190 -611 -185
rect -634 -191 -614 -190
rect -638 -192 -614 -191
rect -612 -192 -611 -190
rect -638 -194 -611 -192
rect -606 -190 -600 -189
rect -606 -192 -604 -190
rect -602 -192 -600 -190
rect -606 -200 -600 -192
rect -584 -182 -578 -181
rect -584 -184 -582 -182
rect -580 -184 -578 -182
rect -584 -189 -578 -184
rect -556 -181 -552 -178
rect -561 -183 -552 -181
rect -541 -182 -540 -176
rect -494 -153 -490 -144
rect -453 -150 -423 -149
rect -453 -152 -451 -150
rect -449 -152 -423 -150
rect -453 -153 -423 -152
rect -494 -155 -493 -153
rect -491 -155 -490 -153
rect -494 -157 -490 -155
rect -427 -157 -423 -153
rect -561 -185 -560 -183
rect -558 -185 -552 -183
rect -427 -161 -418 -157
rect -415 -161 -414 -155
rect -404 -155 -400 -144
rect -404 -157 -403 -155
rect -401 -157 -400 -155
rect -404 -159 -400 -157
rect -422 -167 -418 -161
rect -422 -169 -421 -167
rect -419 -169 -418 -167
rect -443 -174 -437 -173
rect -422 -174 -418 -169
rect -430 -178 -418 -174
rect -584 -191 -582 -189
rect -580 -190 -578 -189
rect -561 -190 -557 -185
rect -580 -191 -560 -190
rect -584 -192 -560 -191
rect -558 -192 -557 -190
rect -584 -194 -557 -192
rect -552 -190 -546 -189
rect -552 -192 -550 -190
rect -548 -192 -546 -190
rect -552 -200 -546 -192
rect -458 -182 -452 -181
rect -458 -184 -456 -182
rect -454 -184 -452 -182
rect -529 -191 -525 -189
rect -529 -193 -528 -191
rect -526 -193 -525 -191
rect -529 -198 -525 -193
rect -494 -191 -490 -189
rect -494 -193 -493 -191
rect -491 -193 -490 -191
rect -529 -200 -528 -198
rect -526 -200 -525 -198
rect -494 -198 -490 -193
rect -458 -189 -452 -184
rect -430 -181 -426 -178
rect -435 -183 -426 -181
rect -415 -182 -414 -176
rect -390 -162 -389 -156
rect -378 -155 -374 -144
rect -378 -157 -377 -155
rect -375 -157 -374 -155
rect -378 -159 -374 -157
rect -364 -162 -363 -156
rect -348 -150 -318 -149
rect -348 -152 -346 -150
rect -344 -152 -318 -150
rect -348 -153 -318 -152
rect -322 -157 -318 -153
rect -390 -181 -389 -174
rect -364 -181 -363 -174
rect -322 -161 -313 -157
rect -310 -161 -309 -155
rect -294 -150 -264 -149
rect -294 -152 -292 -150
rect -290 -152 -264 -150
rect -294 -153 -264 -152
rect -268 -157 -264 -153
rect -317 -167 -313 -161
rect -317 -169 -316 -167
rect -314 -169 -313 -167
rect -338 -174 -332 -173
rect -317 -174 -313 -169
rect -325 -178 -313 -174
rect -435 -185 -434 -183
rect -432 -185 -426 -183
rect -458 -191 -456 -189
rect -454 -190 -452 -189
rect -435 -190 -431 -185
rect -353 -182 -347 -181
rect -353 -184 -351 -182
rect -349 -184 -347 -182
rect -454 -191 -434 -190
rect -458 -192 -434 -191
rect -432 -192 -431 -190
rect -458 -194 -431 -192
rect -426 -190 -420 -189
rect -426 -192 -424 -190
rect -422 -192 -420 -190
rect -494 -200 -493 -198
rect -491 -200 -490 -198
rect -426 -200 -420 -192
rect -353 -189 -347 -184
rect -325 -181 -321 -178
rect -330 -183 -321 -181
rect -310 -182 -309 -176
rect -268 -161 -259 -157
rect -256 -161 -255 -155
rect -244 -153 -240 -144
rect -244 -155 -243 -153
rect -241 -155 -240 -153
rect -244 -157 -240 -155
rect -263 -167 -259 -161
rect -263 -169 -262 -167
rect -260 -169 -259 -167
rect -284 -174 -278 -173
rect -263 -174 -259 -169
rect -271 -178 -259 -174
rect -330 -185 -329 -183
rect -327 -185 -321 -183
rect -402 -191 -396 -190
rect -402 -193 -400 -191
rect -398 -193 -396 -191
rect -402 -200 -396 -193
rect -376 -191 -370 -190
rect -376 -193 -374 -191
rect -372 -193 -370 -191
rect -376 -200 -370 -193
rect -353 -191 -351 -189
rect -349 -190 -347 -189
rect -330 -190 -326 -185
rect -349 -191 -329 -190
rect -353 -192 -329 -191
rect -327 -192 -326 -190
rect -353 -194 -326 -192
rect -321 -190 -315 -189
rect -321 -192 -319 -190
rect -317 -192 -315 -190
rect -321 -200 -315 -192
rect -299 -182 -293 -181
rect -299 -184 -297 -182
rect -295 -184 -293 -182
rect -299 -189 -293 -184
rect -271 -181 -267 -178
rect -276 -183 -267 -181
rect -256 -182 -255 -176
rect -209 -153 -205 -144
rect -168 -150 -138 -149
rect -168 -152 -166 -150
rect -164 -152 -138 -150
rect -168 -153 -138 -152
rect -209 -155 -208 -153
rect -206 -155 -205 -153
rect -209 -157 -205 -155
rect -142 -157 -138 -153
rect -276 -185 -275 -183
rect -273 -185 -267 -183
rect -142 -161 -133 -157
rect -130 -161 -129 -155
rect -119 -155 -115 -144
rect -119 -157 -118 -155
rect -116 -157 -115 -155
rect -119 -159 -115 -157
rect -137 -167 -133 -161
rect -137 -169 -136 -167
rect -134 -169 -133 -167
rect -158 -174 -152 -173
rect -137 -174 -133 -169
rect -145 -178 -133 -174
rect -299 -191 -297 -189
rect -295 -190 -293 -189
rect -276 -190 -272 -185
rect -295 -191 -275 -190
rect -299 -192 -275 -191
rect -273 -192 -272 -190
rect -299 -194 -272 -192
rect -267 -190 -261 -189
rect -267 -192 -265 -190
rect -263 -192 -261 -190
rect -267 -200 -261 -192
rect -173 -182 -167 -181
rect -173 -184 -171 -182
rect -169 -184 -167 -182
rect -244 -191 -240 -189
rect -244 -193 -243 -191
rect -241 -193 -240 -191
rect -244 -198 -240 -193
rect -209 -191 -205 -189
rect -209 -193 -208 -191
rect -206 -193 -205 -191
rect -244 -200 -243 -198
rect -241 -200 -240 -198
rect -209 -198 -205 -193
rect -173 -189 -167 -184
rect -145 -181 -141 -178
rect -150 -183 -141 -181
rect -130 -182 -129 -176
rect -105 -162 -104 -156
rect -93 -155 -89 -144
rect -93 -157 -92 -155
rect -90 -157 -89 -155
rect -93 -159 -89 -157
rect -79 -162 -78 -156
rect -63 -150 -33 -149
rect -63 -152 -61 -150
rect -59 -152 -33 -150
rect -63 -153 -33 -152
rect -37 -157 -33 -153
rect -105 -181 -104 -174
rect -79 -181 -78 -174
rect -37 -161 -28 -157
rect -25 -161 -24 -155
rect -9 -150 21 -149
rect -9 -152 -7 -150
rect -5 -152 21 -150
rect -9 -153 21 -152
rect 17 -157 21 -153
rect -32 -167 -28 -161
rect -32 -169 -31 -167
rect -29 -169 -28 -167
rect -53 -174 -47 -173
rect -32 -174 -28 -169
rect -40 -178 -28 -174
rect -150 -185 -149 -183
rect -147 -185 -141 -183
rect -173 -191 -171 -189
rect -169 -190 -167 -189
rect -150 -190 -146 -185
rect -68 -182 -62 -181
rect -68 -184 -66 -182
rect -64 -184 -62 -182
rect -169 -191 -149 -190
rect -173 -192 -149 -191
rect -147 -192 -146 -190
rect -173 -194 -146 -192
rect -141 -190 -135 -189
rect -141 -192 -139 -190
rect -137 -192 -135 -190
rect -209 -200 -208 -198
rect -206 -200 -205 -198
rect -141 -200 -135 -192
rect -68 -189 -62 -184
rect -40 -181 -36 -178
rect -45 -183 -36 -181
rect -25 -182 -24 -176
rect 17 -161 26 -157
rect 29 -161 30 -155
rect 41 -153 45 -144
rect 41 -155 42 -153
rect 44 -155 45 -153
rect 41 -157 45 -155
rect 22 -167 26 -161
rect 22 -169 23 -167
rect 25 -169 26 -167
rect 1 -174 7 -173
rect 22 -174 26 -169
rect 14 -178 26 -174
rect -45 -185 -44 -183
rect -42 -185 -36 -183
rect -117 -191 -111 -190
rect -117 -193 -115 -191
rect -113 -193 -111 -191
rect -117 -200 -111 -193
rect -91 -191 -85 -190
rect -91 -193 -89 -191
rect -87 -193 -85 -191
rect -91 -200 -85 -193
rect -68 -191 -66 -189
rect -64 -190 -62 -189
rect -45 -190 -41 -185
rect -64 -191 -44 -190
rect -68 -192 -44 -191
rect -42 -192 -41 -190
rect -68 -194 -41 -192
rect -36 -190 -30 -189
rect -36 -192 -34 -190
rect -32 -192 -30 -190
rect -36 -200 -30 -192
rect -14 -182 -8 -181
rect -14 -184 -12 -182
rect -10 -184 -8 -182
rect -14 -189 -8 -184
rect 14 -181 18 -178
rect 9 -183 18 -181
rect 29 -182 30 -176
rect 76 -153 80 -144
rect 117 -150 147 -149
rect 117 -152 119 -150
rect 121 -152 147 -150
rect 117 -153 147 -152
rect 76 -155 77 -153
rect 79 -155 80 -153
rect 76 -157 80 -155
rect 143 -157 147 -153
rect 9 -185 10 -183
rect 12 -185 18 -183
rect 143 -161 152 -157
rect 155 -161 156 -155
rect 166 -155 170 -144
rect 166 -157 167 -155
rect 169 -157 170 -155
rect 166 -159 170 -157
rect 148 -167 152 -161
rect 148 -169 149 -167
rect 151 -169 152 -167
rect 127 -174 133 -173
rect 148 -174 152 -169
rect 140 -178 152 -174
rect -14 -191 -12 -189
rect -10 -190 -8 -189
rect 9 -190 13 -185
rect -10 -191 10 -190
rect -14 -192 10 -191
rect 12 -192 13 -190
rect -14 -194 13 -192
rect 18 -190 24 -189
rect 18 -192 20 -190
rect 22 -192 24 -190
rect 18 -200 24 -192
rect 112 -182 118 -181
rect 112 -184 114 -182
rect 116 -184 118 -182
rect 41 -191 45 -189
rect 41 -193 42 -191
rect 44 -193 45 -191
rect 41 -198 45 -193
rect 76 -191 80 -189
rect 76 -193 77 -191
rect 79 -193 80 -191
rect 41 -200 42 -198
rect 44 -200 45 -198
rect 76 -198 80 -193
rect 112 -189 118 -184
rect 140 -181 144 -178
rect 135 -183 144 -181
rect 155 -182 156 -176
rect 180 -162 181 -156
rect 192 -155 196 -144
rect 192 -157 193 -155
rect 195 -157 196 -155
rect 192 -159 196 -157
rect 206 -162 207 -156
rect 222 -150 252 -149
rect 222 -152 224 -150
rect 226 -152 252 -150
rect 222 -153 252 -152
rect 248 -157 252 -153
rect 180 -181 181 -174
rect 206 -181 207 -174
rect 248 -161 257 -157
rect 260 -161 261 -155
rect 276 -150 306 -149
rect 276 -152 278 -150
rect 280 -152 306 -150
rect 276 -153 306 -152
rect 302 -157 306 -153
rect 253 -167 257 -161
rect 253 -169 254 -167
rect 256 -169 257 -167
rect 232 -174 238 -173
rect 253 -174 257 -169
rect 245 -178 257 -174
rect 135 -185 136 -183
rect 138 -185 144 -183
rect 112 -191 114 -189
rect 116 -190 118 -189
rect 135 -190 139 -185
rect 217 -182 223 -181
rect 217 -184 219 -182
rect 221 -184 223 -182
rect 116 -191 136 -190
rect 112 -192 136 -191
rect 138 -192 139 -190
rect 112 -194 139 -192
rect 144 -190 150 -189
rect 144 -192 146 -190
rect 148 -192 150 -190
rect 76 -200 77 -198
rect 79 -200 80 -198
rect 144 -200 150 -192
rect 217 -189 223 -184
rect 245 -181 249 -178
rect 240 -183 249 -181
rect 260 -182 261 -176
rect 302 -161 311 -157
rect 314 -161 315 -155
rect 326 -153 330 -144
rect 326 -155 327 -153
rect 329 -155 330 -153
rect 326 -157 330 -155
rect 307 -167 311 -161
rect 307 -169 308 -167
rect 310 -169 311 -167
rect 286 -174 292 -173
rect 307 -174 311 -169
rect 299 -178 311 -174
rect 240 -185 241 -183
rect 243 -185 249 -183
rect 168 -191 174 -190
rect 168 -193 170 -191
rect 172 -193 174 -191
rect 168 -200 174 -193
rect 194 -191 200 -190
rect 194 -193 196 -191
rect 198 -193 200 -191
rect 194 -200 200 -193
rect 217 -191 219 -189
rect 221 -190 223 -189
rect 240 -190 244 -185
rect 221 -191 241 -190
rect 217 -192 241 -191
rect 243 -192 244 -190
rect 217 -194 244 -192
rect 249 -190 255 -189
rect 249 -192 251 -190
rect 253 -192 255 -190
rect 249 -200 255 -192
rect 271 -182 277 -181
rect 271 -184 273 -182
rect 275 -184 277 -182
rect 271 -189 277 -184
rect 299 -181 303 -178
rect 294 -183 303 -181
rect 314 -182 315 -176
rect 361 -153 365 -144
rect 402 -150 432 -149
rect 402 -152 404 -150
rect 406 -152 432 -150
rect 402 -153 432 -152
rect 361 -155 362 -153
rect 364 -155 365 -153
rect 361 -157 365 -155
rect 428 -157 432 -153
rect 294 -185 295 -183
rect 297 -185 303 -183
rect 428 -161 437 -157
rect 440 -161 441 -155
rect 488 -150 521 -149
rect 488 -152 490 -150
rect 492 -152 512 -150
rect 514 -152 521 -150
rect 488 -153 521 -152
rect 433 -167 437 -161
rect 433 -169 434 -167
rect 436 -169 437 -167
rect 412 -174 418 -173
rect 433 -174 437 -169
rect 425 -178 437 -174
rect 271 -191 273 -189
rect 275 -190 277 -189
rect 294 -190 298 -185
rect 275 -191 295 -190
rect 271 -192 295 -191
rect 297 -192 298 -190
rect 271 -194 298 -192
rect 303 -190 309 -189
rect 303 -192 305 -190
rect 307 -192 309 -190
rect 303 -200 309 -192
rect 397 -182 403 -181
rect 397 -184 399 -182
rect 401 -184 403 -182
rect 326 -191 330 -189
rect 326 -193 327 -191
rect 329 -193 330 -191
rect 326 -198 330 -193
rect 361 -191 365 -189
rect 361 -193 362 -191
rect 364 -193 365 -191
rect 326 -200 327 -198
rect 329 -200 330 -198
rect 361 -198 365 -193
rect 397 -189 403 -184
rect 425 -181 429 -178
rect 420 -183 429 -181
rect 440 -182 441 -176
rect 517 -160 521 -153
rect 517 -162 530 -160
rect 517 -164 527 -162
rect 529 -164 530 -162
rect 420 -185 421 -183
rect 423 -185 429 -183
rect 397 -191 399 -189
rect 401 -190 403 -189
rect 420 -190 424 -185
rect 517 -182 518 -171
rect 401 -191 421 -190
rect 397 -192 421 -191
rect 423 -192 424 -190
rect 397 -194 424 -192
rect 429 -190 435 -189
rect 429 -192 431 -190
rect 433 -192 435 -190
rect 361 -200 362 -198
rect 364 -200 365 -198
rect 429 -200 435 -192
rect 459 -196 463 -194
rect 526 -190 530 -164
rect 580 -150 613 -149
rect 580 -152 582 -150
rect 584 -152 604 -150
rect 606 -152 613 -150
rect 580 -153 613 -152
rect 533 -187 534 -174
rect 609 -160 613 -153
rect 609 -162 622 -160
rect 609 -164 619 -162
rect 621 -164 622 -162
rect 489 -191 530 -190
rect 489 -193 491 -191
rect 493 -193 530 -191
rect 489 -194 530 -193
rect 609 -182 610 -171
rect 459 -198 460 -196
rect 462 -198 463 -196
rect 551 -196 555 -194
rect 618 -190 622 -164
rect 625 -187 626 -174
rect 581 -191 622 -190
rect 581 -193 583 -191
rect 585 -193 622 -191
rect 581 -194 622 -193
rect 459 -200 463 -198
rect 521 -198 527 -197
rect 521 -200 523 -198
rect 525 -200 527 -198
rect 551 -198 552 -196
rect 554 -198 555 -196
rect 551 -200 555 -198
rect 613 -198 619 -197
rect 613 -200 615 -198
rect 617 -200 619 -198
rect -687 -223 -681 -216
rect -687 -225 -685 -223
rect -683 -225 -681 -223
rect -687 -226 -681 -225
rect -661 -223 -655 -216
rect -661 -225 -659 -223
rect -657 -225 -655 -223
rect -661 -226 -655 -225
rect -638 -224 -611 -222
rect -638 -225 -614 -224
rect -638 -227 -636 -225
rect -634 -226 -614 -225
rect -612 -226 -611 -224
rect -634 -227 -632 -226
rect -638 -232 -632 -227
rect -638 -234 -636 -232
rect -634 -234 -632 -232
rect -638 -235 -632 -234
rect -675 -242 -674 -235
rect -689 -259 -685 -257
rect -649 -242 -648 -235
rect -615 -231 -611 -226
rect -606 -224 -600 -216
rect -606 -226 -604 -224
rect -602 -226 -600 -224
rect -606 -227 -600 -226
rect -615 -233 -614 -231
rect -612 -233 -606 -231
rect -615 -235 -606 -233
rect -610 -238 -606 -235
rect -689 -261 -688 -259
rect -686 -261 -685 -259
rect -675 -260 -674 -254
rect -689 -272 -685 -261
rect -663 -259 -659 -257
rect -610 -242 -598 -238
rect -595 -240 -594 -234
rect -584 -224 -557 -222
rect -584 -225 -560 -224
rect -584 -227 -582 -225
rect -580 -226 -560 -225
rect -558 -226 -557 -224
rect -580 -227 -578 -226
rect -584 -232 -578 -227
rect -584 -234 -582 -232
rect -580 -234 -578 -232
rect -584 -235 -578 -234
rect -561 -231 -557 -226
rect -552 -224 -546 -216
rect -529 -218 -528 -216
rect -526 -218 -525 -216
rect -552 -226 -550 -224
rect -548 -226 -546 -224
rect -552 -227 -546 -226
rect -529 -223 -525 -218
rect -494 -218 -493 -216
rect -491 -218 -490 -216
rect -529 -225 -528 -223
rect -526 -225 -525 -223
rect -529 -227 -525 -225
rect -561 -233 -560 -231
rect -558 -233 -552 -231
rect -561 -235 -552 -233
rect -494 -223 -490 -218
rect -494 -225 -493 -223
rect -491 -225 -490 -223
rect -494 -227 -490 -225
rect -458 -224 -431 -222
rect -458 -225 -434 -224
rect -458 -227 -456 -225
rect -454 -226 -434 -225
rect -432 -226 -431 -224
rect -454 -227 -452 -226
rect -556 -238 -552 -235
rect -623 -243 -617 -242
rect -663 -261 -662 -259
rect -660 -261 -659 -259
rect -649 -260 -648 -254
rect -663 -272 -659 -261
rect -602 -247 -598 -242
rect -602 -249 -601 -247
rect -599 -249 -598 -247
rect -602 -255 -598 -249
rect -556 -242 -544 -238
rect -541 -240 -540 -234
rect -569 -243 -563 -242
rect -607 -259 -598 -255
rect -607 -263 -603 -259
rect -595 -261 -594 -255
rect -548 -247 -544 -242
rect -548 -249 -547 -247
rect -545 -249 -544 -247
rect -548 -255 -544 -249
rect -553 -259 -544 -255
rect -633 -264 -603 -263
rect -633 -266 -631 -264
rect -629 -266 -603 -264
rect -633 -267 -603 -266
rect -553 -263 -549 -259
rect -541 -261 -540 -255
rect -579 -264 -549 -263
rect -579 -266 -577 -264
rect -575 -266 -549 -264
rect -579 -267 -549 -266
rect -529 -261 -525 -259
rect -458 -232 -452 -227
rect -458 -234 -456 -232
rect -454 -234 -452 -232
rect -458 -235 -452 -234
rect -435 -231 -431 -226
rect -426 -224 -420 -216
rect -426 -226 -424 -224
rect -422 -226 -420 -224
rect -426 -227 -420 -226
rect -402 -223 -396 -216
rect -402 -225 -400 -223
rect -398 -225 -396 -223
rect -402 -226 -396 -225
rect -376 -223 -370 -216
rect -376 -225 -374 -223
rect -372 -225 -370 -223
rect -376 -226 -370 -225
rect -353 -224 -326 -222
rect -353 -225 -329 -224
rect -353 -227 -351 -225
rect -349 -226 -329 -225
rect -327 -226 -326 -224
rect -349 -227 -347 -226
rect -435 -233 -434 -231
rect -432 -233 -426 -231
rect -435 -235 -426 -233
rect -430 -238 -426 -235
rect -430 -242 -418 -238
rect -415 -240 -414 -234
rect -353 -232 -347 -227
rect -353 -234 -351 -232
rect -349 -234 -347 -232
rect -353 -235 -347 -234
rect -443 -243 -437 -242
rect -422 -247 -418 -242
rect -422 -249 -421 -247
rect -419 -249 -418 -247
rect -422 -255 -418 -249
rect -390 -242 -389 -235
rect -427 -259 -418 -255
rect -529 -263 -528 -261
rect -526 -263 -525 -261
rect -529 -272 -525 -263
rect -494 -261 -490 -259
rect -494 -263 -493 -261
rect -491 -263 -490 -261
rect -427 -263 -423 -259
rect -415 -261 -414 -255
rect -494 -272 -490 -263
rect -453 -264 -423 -263
rect -453 -266 -451 -264
rect -449 -266 -423 -264
rect -453 -267 -423 -266
rect -404 -259 -400 -257
rect -364 -242 -363 -235
rect -330 -231 -326 -226
rect -321 -224 -315 -216
rect -321 -226 -319 -224
rect -317 -226 -315 -224
rect -321 -227 -315 -226
rect -330 -233 -329 -231
rect -327 -233 -321 -231
rect -330 -235 -321 -233
rect -325 -238 -321 -235
rect -404 -261 -403 -259
rect -401 -261 -400 -259
rect -390 -260 -389 -254
rect -404 -272 -400 -261
rect -378 -259 -374 -257
rect -325 -242 -313 -238
rect -310 -240 -309 -234
rect -299 -224 -272 -222
rect -299 -225 -275 -224
rect -299 -227 -297 -225
rect -295 -226 -275 -225
rect -273 -226 -272 -224
rect -295 -227 -293 -226
rect -299 -232 -293 -227
rect -299 -234 -297 -232
rect -295 -234 -293 -232
rect -299 -235 -293 -234
rect -276 -231 -272 -226
rect -267 -224 -261 -216
rect -244 -218 -243 -216
rect -241 -218 -240 -216
rect -267 -226 -265 -224
rect -263 -226 -261 -224
rect -267 -227 -261 -226
rect -244 -223 -240 -218
rect -209 -218 -208 -216
rect -206 -218 -205 -216
rect -244 -225 -243 -223
rect -241 -225 -240 -223
rect -244 -227 -240 -225
rect -276 -233 -275 -231
rect -273 -233 -267 -231
rect -276 -235 -267 -233
rect -209 -223 -205 -218
rect -209 -225 -208 -223
rect -206 -225 -205 -223
rect -209 -227 -205 -225
rect -173 -224 -146 -222
rect -173 -225 -149 -224
rect -173 -227 -171 -225
rect -169 -226 -149 -225
rect -147 -226 -146 -224
rect -169 -227 -167 -226
rect -271 -238 -267 -235
rect -338 -243 -332 -242
rect -378 -261 -377 -259
rect -375 -261 -374 -259
rect -364 -260 -363 -254
rect -378 -272 -374 -261
rect -317 -247 -313 -242
rect -317 -249 -316 -247
rect -314 -249 -313 -247
rect -317 -255 -313 -249
rect -271 -242 -259 -238
rect -256 -240 -255 -234
rect -284 -243 -278 -242
rect -322 -259 -313 -255
rect -322 -263 -318 -259
rect -310 -261 -309 -255
rect -263 -247 -259 -242
rect -263 -249 -262 -247
rect -260 -249 -259 -247
rect -263 -255 -259 -249
rect -268 -259 -259 -255
rect -348 -264 -318 -263
rect -348 -266 -346 -264
rect -344 -266 -318 -264
rect -348 -267 -318 -266
rect -268 -263 -264 -259
rect -256 -261 -255 -255
rect -294 -264 -264 -263
rect -294 -266 -292 -264
rect -290 -266 -264 -264
rect -294 -267 -264 -266
rect -244 -261 -240 -259
rect -173 -232 -167 -227
rect -173 -234 -171 -232
rect -169 -234 -167 -232
rect -173 -235 -167 -234
rect -150 -231 -146 -226
rect -141 -224 -135 -216
rect -141 -226 -139 -224
rect -137 -226 -135 -224
rect -141 -227 -135 -226
rect -117 -223 -111 -216
rect -117 -225 -115 -223
rect -113 -225 -111 -223
rect -117 -226 -111 -225
rect -91 -223 -85 -216
rect -91 -225 -89 -223
rect -87 -225 -85 -223
rect -91 -226 -85 -225
rect -68 -224 -41 -222
rect -68 -225 -44 -224
rect -68 -227 -66 -225
rect -64 -226 -44 -225
rect -42 -226 -41 -224
rect -64 -227 -62 -226
rect -150 -233 -149 -231
rect -147 -233 -141 -231
rect -150 -235 -141 -233
rect -145 -238 -141 -235
rect -145 -242 -133 -238
rect -130 -240 -129 -234
rect -68 -232 -62 -227
rect -68 -234 -66 -232
rect -64 -234 -62 -232
rect -68 -235 -62 -234
rect -158 -243 -152 -242
rect -137 -247 -133 -242
rect -137 -249 -136 -247
rect -134 -249 -133 -247
rect -137 -255 -133 -249
rect -105 -242 -104 -235
rect -142 -259 -133 -255
rect -244 -263 -243 -261
rect -241 -263 -240 -261
rect -244 -272 -240 -263
rect -209 -261 -205 -259
rect -209 -263 -208 -261
rect -206 -263 -205 -261
rect -142 -263 -138 -259
rect -130 -261 -129 -255
rect -209 -272 -205 -263
rect -168 -264 -138 -263
rect -168 -266 -166 -264
rect -164 -266 -138 -264
rect -168 -267 -138 -266
rect -119 -259 -115 -257
rect -79 -242 -78 -235
rect -45 -231 -41 -226
rect -36 -224 -30 -216
rect -36 -226 -34 -224
rect -32 -226 -30 -224
rect -36 -227 -30 -226
rect -45 -233 -44 -231
rect -42 -233 -36 -231
rect -45 -235 -36 -233
rect -40 -238 -36 -235
rect -119 -261 -118 -259
rect -116 -261 -115 -259
rect -105 -260 -104 -254
rect -119 -272 -115 -261
rect -93 -259 -89 -257
rect -40 -242 -28 -238
rect -25 -240 -24 -234
rect -14 -224 13 -222
rect -14 -225 10 -224
rect -14 -227 -12 -225
rect -10 -226 10 -225
rect 12 -226 13 -224
rect -10 -227 -8 -226
rect -14 -232 -8 -227
rect -14 -234 -12 -232
rect -10 -234 -8 -232
rect -14 -235 -8 -234
rect 9 -231 13 -226
rect 18 -224 24 -216
rect 41 -218 42 -216
rect 44 -218 45 -216
rect 18 -226 20 -224
rect 22 -226 24 -224
rect 18 -227 24 -226
rect 41 -223 45 -218
rect 76 -218 77 -216
rect 79 -218 80 -216
rect 41 -225 42 -223
rect 44 -225 45 -223
rect 41 -227 45 -225
rect 9 -233 10 -231
rect 12 -233 18 -231
rect 9 -235 18 -233
rect 76 -223 80 -218
rect 76 -225 77 -223
rect 79 -225 80 -223
rect 76 -227 80 -225
rect 112 -224 139 -222
rect 112 -225 136 -224
rect 112 -227 114 -225
rect 116 -226 136 -225
rect 138 -226 139 -224
rect 116 -227 118 -226
rect 14 -238 18 -235
rect -53 -243 -47 -242
rect -93 -261 -92 -259
rect -90 -261 -89 -259
rect -79 -260 -78 -254
rect -93 -272 -89 -261
rect -32 -247 -28 -242
rect -32 -249 -31 -247
rect -29 -249 -28 -247
rect -32 -255 -28 -249
rect 14 -242 26 -238
rect 29 -240 30 -234
rect 1 -243 7 -242
rect -37 -259 -28 -255
rect -37 -263 -33 -259
rect -25 -261 -24 -255
rect 22 -247 26 -242
rect 22 -249 23 -247
rect 25 -249 26 -247
rect 22 -255 26 -249
rect 17 -259 26 -255
rect -63 -264 -33 -263
rect -63 -266 -61 -264
rect -59 -266 -33 -264
rect -63 -267 -33 -266
rect 17 -263 21 -259
rect 29 -261 30 -255
rect -9 -264 21 -263
rect -9 -266 -7 -264
rect -5 -266 21 -264
rect -9 -267 21 -266
rect 41 -261 45 -259
rect 112 -232 118 -227
rect 112 -234 114 -232
rect 116 -234 118 -232
rect 112 -235 118 -234
rect 135 -231 139 -226
rect 144 -224 150 -216
rect 144 -226 146 -224
rect 148 -226 150 -224
rect 144 -227 150 -226
rect 168 -223 174 -216
rect 168 -225 170 -223
rect 172 -225 174 -223
rect 168 -226 174 -225
rect 194 -223 200 -216
rect 194 -225 196 -223
rect 198 -225 200 -223
rect 194 -226 200 -225
rect 217 -224 244 -222
rect 217 -225 241 -224
rect 217 -227 219 -225
rect 221 -226 241 -225
rect 243 -226 244 -224
rect 221 -227 223 -226
rect 135 -233 136 -231
rect 138 -233 144 -231
rect 135 -235 144 -233
rect 140 -238 144 -235
rect 140 -242 152 -238
rect 155 -240 156 -234
rect 217 -232 223 -227
rect 217 -234 219 -232
rect 221 -234 223 -232
rect 217 -235 223 -234
rect 127 -243 133 -242
rect 148 -247 152 -242
rect 148 -249 149 -247
rect 151 -249 152 -247
rect 148 -255 152 -249
rect 180 -242 181 -235
rect 143 -259 152 -255
rect 41 -263 42 -261
rect 44 -263 45 -261
rect 41 -272 45 -263
rect 76 -261 80 -259
rect 76 -263 77 -261
rect 79 -263 80 -261
rect 143 -263 147 -259
rect 155 -261 156 -255
rect 76 -272 80 -263
rect 117 -264 147 -263
rect 117 -266 119 -264
rect 121 -266 147 -264
rect 117 -267 147 -266
rect 166 -259 170 -257
rect 206 -242 207 -235
rect 240 -231 244 -226
rect 249 -224 255 -216
rect 249 -226 251 -224
rect 253 -226 255 -224
rect 249 -227 255 -226
rect 240 -233 241 -231
rect 243 -233 249 -231
rect 240 -235 249 -233
rect 245 -238 249 -235
rect 166 -261 167 -259
rect 169 -261 170 -259
rect 180 -260 181 -254
rect 166 -272 170 -261
rect 192 -259 196 -257
rect 245 -242 257 -238
rect 260 -240 261 -234
rect 271 -224 298 -222
rect 271 -225 295 -224
rect 271 -227 273 -225
rect 275 -226 295 -225
rect 297 -226 298 -224
rect 275 -227 277 -226
rect 271 -232 277 -227
rect 271 -234 273 -232
rect 275 -234 277 -232
rect 271 -235 277 -234
rect 294 -231 298 -226
rect 303 -224 309 -216
rect 326 -218 327 -216
rect 329 -218 330 -216
rect 303 -226 305 -224
rect 307 -226 309 -224
rect 303 -227 309 -226
rect 326 -223 330 -218
rect 361 -218 362 -216
rect 364 -218 365 -216
rect 326 -225 327 -223
rect 329 -225 330 -223
rect 326 -227 330 -225
rect 294 -233 295 -231
rect 297 -233 303 -231
rect 294 -235 303 -233
rect 361 -223 365 -218
rect 361 -225 362 -223
rect 364 -225 365 -223
rect 361 -227 365 -225
rect 397 -224 424 -222
rect 397 -225 421 -224
rect 397 -227 399 -225
rect 401 -226 421 -225
rect 423 -226 424 -224
rect 401 -227 403 -226
rect 299 -238 303 -235
rect 232 -243 238 -242
rect 192 -261 193 -259
rect 195 -261 196 -259
rect 206 -260 207 -254
rect 192 -272 196 -261
rect 253 -247 257 -242
rect 253 -249 254 -247
rect 256 -249 257 -247
rect 253 -255 257 -249
rect 299 -242 311 -238
rect 314 -240 315 -234
rect 286 -243 292 -242
rect 248 -259 257 -255
rect 248 -263 252 -259
rect 260 -261 261 -255
rect 307 -247 311 -242
rect 307 -249 308 -247
rect 310 -249 311 -247
rect 307 -255 311 -249
rect 302 -259 311 -255
rect 222 -264 252 -263
rect 222 -266 224 -264
rect 226 -266 252 -264
rect 222 -267 252 -266
rect 302 -263 306 -259
rect 314 -261 315 -255
rect 276 -264 306 -263
rect 276 -266 278 -264
rect 280 -266 306 -264
rect 276 -267 306 -266
rect 326 -261 330 -259
rect 397 -232 403 -227
rect 397 -234 399 -232
rect 401 -234 403 -232
rect 397 -235 403 -234
rect 420 -231 424 -226
rect 429 -224 435 -216
rect 459 -218 463 -216
rect 459 -220 460 -218
rect 462 -220 463 -218
rect 521 -218 523 -216
rect 525 -218 527 -216
rect 521 -219 527 -218
rect 551 -218 555 -216
rect 429 -226 431 -224
rect 433 -226 435 -224
rect 429 -227 435 -226
rect 459 -222 463 -220
rect 551 -220 552 -218
rect 554 -220 555 -218
rect 613 -218 615 -216
rect 617 -218 619 -216
rect 613 -219 619 -218
rect 489 -223 530 -222
rect 489 -225 491 -223
rect 493 -225 530 -223
rect 489 -226 530 -225
rect 420 -233 421 -231
rect 423 -233 429 -231
rect 420 -235 429 -233
rect 425 -238 429 -235
rect 425 -242 437 -238
rect 440 -240 441 -234
rect 412 -243 418 -242
rect 433 -247 437 -242
rect 433 -249 434 -247
rect 436 -249 437 -247
rect 433 -255 437 -249
rect 517 -245 518 -234
rect 526 -252 530 -226
rect 533 -242 534 -229
rect 551 -222 555 -220
rect 581 -223 622 -222
rect 581 -225 583 -223
rect 585 -225 622 -223
rect 581 -226 622 -225
rect 428 -259 437 -255
rect 326 -263 327 -261
rect 329 -263 330 -261
rect 326 -272 330 -263
rect 361 -261 365 -259
rect 361 -263 362 -261
rect 364 -263 365 -261
rect 428 -263 432 -259
rect 440 -261 441 -255
rect 361 -272 365 -263
rect 402 -264 432 -263
rect 402 -266 404 -264
rect 406 -266 432 -264
rect 402 -267 432 -266
rect 517 -254 527 -252
rect 529 -254 530 -252
rect 517 -256 530 -254
rect 517 -263 521 -256
rect 609 -245 610 -234
rect 618 -252 622 -226
rect 625 -242 626 -229
rect 488 -264 521 -263
rect 488 -266 490 -264
rect 492 -266 512 -264
rect 514 -266 521 -264
rect 488 -267 521 -266
rect 609 -254 619 -252
rect 621 -254 622 -252
rect 609 -256 622 -254
rect 609 -263 613 -256
rect 580 -264 613 -263
rect 580 -266 582 -264
rect 584 -266 604 -264
rect 606 -266 613 -264
rect 580 -267 613 -266
<< via1 >>
rect 179 316 181 318
rect 673 316 675 318
rect 150 308 152 310
rect 665 308 667 310
rect -103 300 -101 302
rect 150 300 152 302
rect 158 300 160 302
rect 657 300 659 302
rect -714 292 -712 294
rect -688 292 -686 294
rect -413 292 -411 294
rect -126 292 -124 294
rect -118 292 -116 294
rect 649 292 651 294
rect -706 284 -704 286
rect -403 284 -401 286
rect -126 284 -124 286
rect 158 284 160 286
rect 167 284 169 286
rect 641 284 643 286
rect -663 276 -661 278
rect -378 276 -376 278
rect -93 276 -91 278
rect 192 276 194 278
rect 442 276 444 278
rect 681 276 683 278
rect -617 268 -615 270
rect -332 268 -330 270
rect -47 268 -45 270
rect 238 268 240 270
rect 515 268 517 270
rect -617 260 -615 262
rect -563 260 -561 262
rect -437 260 -435 262
rect -332 260 -330 262
rect -278 260 -276 262
rect -152 260 -150 262
rect -47 260 -45 262
rect 7 260 9 262
rect 133 260 135 262
rect 238 260 240 262
rect 292 260 294 262
rect 418 260 420 262
rect 455 260 457 262
rect 633 260 635 262
rect -663 252 -661 254
rect -446 252 -444 254
rect -378 252 -376 254
rect -161 252 -159 254
rect -93 252 -91 254
rect 124 252 126 254
rect 192 252 194 254
rect 409 252 411 254
rect 455 252 457 254
rect 515 252 517 254
rect -593 244 -591 246
rect -482 244 -480 246
rect -308 244 -306 246
rect -197 244 -195 246
rect -23 244 -21 246
rect 88 244 90 246
rect 262 244 264 246
rect 373 244 375 246
rect 479 244 481 246
rect 539 244 541 246
rect 609 244 611 246
rect 157 240 159 242
rect 179 240 181 242
rect -698 236 -696 238
rect -663 236 -661 238
rect -647 236 -645 238
rect -626 236 -624 238
rect -572 236 -570 238
rect -362 236 -360 238
rect -341 236 -339 238
rect -287 236 -285 238
rect -128 236 -126 238
rect -103 236 -101 238
rect -77 236 -75 238
rect -56 236 -54 238
rect -2 236 0 238
rect 208 236 210 238
rect 229 236 231 238
rect 283 236 285 238
rect 551 236 553 238
rect 581 236 583 238
rect 625 236 627 238
rect -688 228 -686 230
rect -580 228 -578 230
rect -513 228 -511 230
rect -470 228 -468 230
rect -454 228 -452 230
rect -403 228 -401 230
rect -295 228 -293 230
rect -228 228 -226 230
rect -185 228 -183 230
rect -169 228 -167 230
rect -118 228 -116 230
rect -10 228 -8 230
rect 57 228 59 230
rect 100 228 102 230
rect 116 228 118 230
rect 167 228 169 230
rect 275 228 277 230
rect 342 228 344 230
rect 385 228 387 230
rect 401 228 403 230
rect 489 228 491 230
rect 597 228 599 230
rect 617 228 619 230
rect -673 220 -671 222
rect -634 220 -632 222
rect -539 220 -537 222
rect -529 220 -527 222
rect -505 220 -503 222
rect -494 220 -492 222
rect -482 220 -480 222
rect -388 220 -386 222
rect -349 220 -347 222
rect -254 220 -252 222
rect -244 220 -242 222
rect -220 220 -218 222
rect -209 220 -207 222
rect -197 220 -195 222
rect -103 220 -101 222
rect -64 220 -62 222
rect 31 220 33 222
rect 41 220 43 222
rect 65 220 67 222
rect 76 220 78 222
rect 88 220 90 222
rect 182 220 184 222
rect 221 220 223 222
rect 316 220 318 222
rect 326 220 328 222
rect 350 220 352 222
rect 361 220 363 222
rect 373 220 375 222
rect 500 220 502 222
rect 560 220 562 222
rect 739 209 741 211
rect -688 181 -686 183
rect -673 184 -671 186
rect -663 181 -661 183
rect -647 184 -645 186
rect -634 190 -632 192
rect -617 188 -615 190
rect -626 173 -624 175
rect -593 183 -591 185
rect -580 190 -578 192
rect -563 188 -561 190
rect -572 173 -570 175
rect -539 183 -537 185
rect -529 184 -527 186
rect -505 189 -503 191
rect -513 176 -511 178
rect -494 184 -492 186
rect -470 191 -468 193
rect -482 176 -480 178
rect -454 190 -452 192
rect -437 189 -435 191
rect -446 173 -444 175
rect -413 187 -411 189
rect -403 181 -401 183
rect -388 184 -386 186
rect -378 181 -376 183
rect -362 184 -360 186
rect -349 190 -347 192
rect -332 188 -330 190
rect -341 173 -339 175
rect -308 183 -306 185
rect -295 190 -293 192
rect -278 188 -276 190
rect -287 173 -285 175
rect -254 183 -252 185
rect -244 184 -242 186
rect -220 189 -218 191
rect -228 176 -226 178
rect -209 184 -207 186
rect -185 191 -183 193
rect -197 176 -195 178
rect -169 190 -167 192
rect -152 189 -150 191
rect -161 173 -159 175
rect -128 187 -126 189
rect -118 181 -116 183
rect -103 184 -101 186
rect -93 181 -91 183
rect -77 184 -75 186
rect -64 190 -62 192
rect -47 188 -45 190
rect -56 173 -54 175
rect -23 183 -21 185
rect -10 190 -8 192
rect 7 188 9 190
rect -2 173 0 175
rect 31 183 33 185
rect 41 184 43 186
rect 65 189 67 191
rect 57 176 59 178
rect 76 184 78 186
rect 100 191 102 193
rect 88 176 90 178
rect 116 190 118 192
rect 133 189 135 191
rect 124 173 126 175
rect 157 187 159 189
rect 167 181 169 183
rect 182 184 184 186
rect 192 181 194 183
rect 208 184 210 186
rect 221 190 223 192
rect 238 188 240 190
rect 229 173 231 175
rect 262 183 264 185
rect 275 190 277 192
rect 292 188 294 190
rect 283 173 285 175
rect 316 183 318 185
rect 326 184 328 186
rect 350 189 352 191
rect 342 176 344 178
rect 361 184 363 186
rect 385 191 387 193
rect 373 176 375 178
rect 401 190 403 192
rect 418 189 420 191
rect 409 173 411 175
rect 442 187 444 189
rect 581 197 583 199
rect 479 190 481 192
rect 455 185 457 187
rect 497 188 499 190
rect 539 190 541 192
rect 515 185 517 187
rect 489 173 491 175
rect 551 190 553 192
rect 560 173 562 175
rect 597 181 599 183
rect -733 141 -731 143
rect -688 101 -686 103
rect -673 98 -671 100
rect -663 101 -661 103
rect -626 109 -624 111
rect -647 98 -645 100
rect -634 92 -632 94
rect -617 94 -615 96
rect -572 109 -570 111
rect -593 99 -591 101
rect -580 92 -578 94
rect -563 94 -561 96
rect -513 106 -511 108
rect -539 99 -537 101
rect -529 98 -527 100
rect -482 106 -480 108
rect -494 98 -492 100
rect -505 93 -503 95
rect -446 109 -444 111
rect -470 91 -468 93
rect -454 92 -452 94
rect -403 101 -401 103
rect -413 95 -411 97
rect -437 93 -435 95
rect -388 98 -386 100
rect -378 101 -376 103
rect -341 109 -339 111
rect -362 98 -360 100
rect -349 92 -347 94
rect -332 94 -330 96
rect -287 109 -285 111
rect -308 99 -306 101
rect -295 92 -293 94
rect -278 94 -276 96
rect -228 106 -226 108
rect -254 99 -252 101
rect -244 98 -242 100
rect -197 106 -195 108
rect -209 98 -207 100
rect -220 93 -218 95
rect -161 109 -159 111
rect -185 91 -183 93
rect -169 92 -167 94
rect -118 101 -116 103
rect -128 95 -126 97
rect -152 93 -150 95
rect -103 98 -101 100
rect -93 101 -91 103
rect -56 109 -54 111
rect -77 98 -75 100
rect -64 92 -62 94
rect -47 94 -45 96
rect -2 109 0 111
rect -23 99 -21 101
rect -10 92 -8 94
rect 7 94 9 96
rect 57 106 59 108
rect 31 99 33 101
rect 41 98 43 100
rect 88 106 90 108
rect 76 98 78 100
rect 65 93 67 95
rect 124 109 126 111
rect 100 91 102 93
rect 116 92 118 94
rect 167 101 169 103
rect 157 95 159 97
rect 133 93 135 95
rect 182 98 184 100
rect 192 101 194 103
rect 229 109 231 111
rect 208 98 210 100
rect 221 92 223 94
rect 238 94 240 96
rect 283 109 285 111
rect 262 99 264 101
rect 275 92 277 94
rect 292 94 294 96
rect 342 106 344 108
rect 316 99 318 101
rect 326 98 328 100
rect 373 106 375 108
rect 361 98 363 100
rect 350 93 352 95
rect 409 109 411 111
rect 385 91 387 93
rect 401 92 403 94
rect 442 95 444 97
rect 418 93 420 95
rect 455 99 457 101
rect 489 109 491 111
rect 515 99 517 101
rect 479 92 481 94
rect 497 94 499 96
rect 549 109 551 111
rect 539 92 541 94
rect 557 94 559 96
rect 597 101 599 103
rect 581 85 583 87
rect 740 73 742 75
rect -673 62 -671 64
rect -634 62 -632 64
rect -539 62 -537 64
rect -529 62 -527 64
rect -505 62 -503 64
rect -494 62 -492 64
rect -482 62 -480 64
rect -388 62 -386 64
rect -349 62 -347 64
rect -254 62 -252 64
rect -244 62 -242 64
rect -220 62 -218 64
rect -209 62 -207 64
rect -197 62 -195 64
rect -103 62 -101 64
rect -64 62 -62 64
rect 31 62 33 64
rect 41 62 43 64
rect 65 62 67 64
rect 76 62 78 64
rect 88 62 90 64
rect 182 62 184 64
rect 221 62 223 64
rect 316 62 318 64
rect 326 62 328 64
rect 350 62 352 64
rect 361 62 363 64
rect 373 62 375 64
rect 500 62 502 64
rect 560 62 562 64
rect -688 54 -686 56
rect -580 54 -578 56
rect -513 54 -511 56
rect -470 54 -468 56
rect -454 54 -452 56
rect -403 54 -401 56
rect -295 54 -293 56
rect -228 54 -226 56
rect -185 54 -183 56
rect -169 54 -167 56
rect -118 54 -116 56
rect -10 54 -8 56
rect 57 54 59 56
rect 100 54 102 56
rect 116 54 118 56
rect 167 54 169 56
rect 275 54 277 56
rect 342 54 344 56
rect 385 54 387 56
rect 401 54 403 56
rect 489 54 491 56
rect 552 54 554 56
rect 597 54 599 56
rect -698 46 -696 48
rect -663 46 -661 48
rect -647 46 -645 48
rect -626 46 -624 48
rect -572 46 -570 48
rect -362 46 -360 48
rect -341 46 -339 48
rect -287 46 -285 48
rect -77 46 -75 48
rect -56 46 -54 48
rect -2 46 0 48
rect 208 46 210 48
rect 229 46 231 48
rect 283 46 285 48
rect 455 46 457 48
rect 515 46 517 48
rect 581 46 583 48
rect 609 46 611 48
rect -593 38 -591 40
rect -482 38 -480 40
rect -308 38 -306 40
rect -197 38 -195 40
rect -23 38 -21 40
rect 88 38 90 40
rect 157 38 159 40
rect 202 38 204 40
rect 262 38 264 40
rect 373 38 375 40
rect 539 38 541 40
rect 617 38 619 40
rect -663 30 -661 32
rect -446 30 -444 32
rect -378 30 -376 32
rect -161 30 -159 32
rect -93 30 -91 32
rect 124 30 126 32
rect 192 30 194 32
rect 409 30 411 32
rect 479 30 481 32
rect 625 30 627 32
rect 681 31 683 33
rect 705 31 707 33
rect -617 22 -615 24
rect -563 22 -561 24
rect -437 22 -435 24
rect -332 22 -330 24
rect -278 22 -276 24
rect -152 22 -150 24
rect -47 22 -45 24
rect 7 22 9 24
rect 133 22 135 24
rect 238 22 240 24
rect 292 22 294 24
rect 418 22 420 24
rect 442 22 444 24
rect 721 22 723 24
rect -617 14 -615 16
rect -332 14 -330 16
rect -47 14 -45 16
rect 238 14 240 16
rect 455 14 457 16
rect -663 6 -661 8
rect -378 6 -376 8
rect -93 6 -91 8
rect 192 6 194 8
rect 202 6 204 8
rect 681 6 683 8
rect -413 -2 -411 0
rect 146 -2 148 0
rect 167 -2 169 0
rect 641 -2 643 0
rect -706 -10 -704 -8
rect -403 -10 -401 -8
rect -128 -10 -126 -8
rect 137 -10 139 -8
rect 146 -10 148 -8
rect 470 -10 472 -8
rect -118 -18 -116 -16
rect 649 -18 651 -16
rect -714 -26 -712 -24
rect -688 -26 -686 -24
rect 137 -26 139 -24
rect 552 -26 554 -24
rect -714 -42 -712 -40
rect -688 -42 -686 -40
rect 157 -42 159 -40
rect 697 -42 699 -40
rect -118 -50 -116 -48
rect 649 -50 651 -48
rect -706 -58 -704 -56
rect -403 -58 -401 -56
rect -128 -58 -126 -56
rect 141 -58 143 -56
rect 149 -58 151 -56
rect 460 -58 462 -56
rect -413 -66 -411 -64
rect 149 -66 151 -64
rect 167 -66 169 -64
rect 641 -66 643 -64
rect -663 -74 -661 -72
rect -378 -74 -376 -72
rect -93 -74 -91 -72
rect 192 -74 194 -72
rect 230 -74 232 -72
rect 562 -74 564 -72
rect -617 -82 -615 -80
rect -332 -82 -330 -80
rect -47 -82 -45 -80
rect 238 -82 240 -80
rect 515 -82 517 -80
rect -617 -90 -615 -88
rect -563 -90 -561 -88
rect -437 -90 -435 -88
rect -332 -90 -330 -88
rect -278 -90 -276 -88
rect -152 -90 -150 -88
rect -47 -90 -45 -88
rect 7 -90 9 -88
rect 133 -90 135 -88
rect 141 -90 143 -88
rect 230 -90 232 -88
rect 238 -90 240 -88
rect 292 -90 294 -88
rect 418 -90 420 -88
rect 442 -90 444 -88
rect 713 -90 715 -88
rect -663 -98 -661 -96
rect -446 -98 -444 -96
rect -378 -98 -376 -96
rect -161 -98 -159 -96
rect -93 -98 -91 -96
rect 124 -98 126 -96
rect 192 -98 194 -96
rect 409 -98 411 -96
rect 681 -98 683 -96
rect 689 -98 691 -96
rect -593 -106 -591 -104
rect -482 -106 -480 -104
rect -308 -106 -306 -104
rect -197 -106 -195 -104
rect -23 -106 -21 -104
rect 88 -106 90 -104
rect 262 -106 264 -104
rect 373 -106 375 -104
rect 591 -106 593 -104
rect 665 -106 667 -104
rect 673 -106 675 -104
rect 681 -106 683 -104
rect -698 -114 -696 -112
rect -663 -114 -661 -112
rect -647 -114 -645 -112
rect -626 -114 -624 -112
rect -572 -114 -570 -112
rect -362 -114 -360 -112
rect -341 -114 -339 -112
rect -287 -114 -285 -112
rect -77 -114 -75 -112
rect -56 -114 -54 -112
rect -2 -114 0 -112
rect 208 -114 210 -112
rect 229 -114 231 -112
rect 283 -114 285 -112
rect 580 -114 582 -112
rect 673 -114 675 -112
rect -688 -122 -686 -120
rect -580 -122 -578 -120
rect -513 -122 -511 -120
rect -470 -122 -468 -120
rect -454 -122 -452 -120
rect -403 -122 -401 -120
rect -295 -122 -293 -120
rect -228 -122 -226 -120
rect -185 -122 -183 -120
rect -169 -122 -167 -120
rect -118 -122 -116 -120
rect -10 -122 -8 -120
rect 57 -122 59 -120
rect 100 -122 102 -120
rect 116 -122 118 -120
rect 167 -122 169 -120
rect 275 -122 277 -120
rect 342 -122 344 -120
rect 385 -122 387 -120
rect 401 -122 403 -120
rect 499 -122 501 -120
rect 665 -122 667 -120
rect -673 -130 -671 -128
rect -634 -130 -632 -128
rect -539 -130 -537 -128
rect -529 -130 -527 -128
rect -505 -130 -503 -128
rect -494 -130 -492 -128
rect -482 -130 -480 -128
rect -388 -130 -386 -128
rect -349 -130 -347 -128
rect -254 -130 -252 -128
rect -244 -130 -242 -128
rect -220 -130 -218 -128
rect -209 -130 -207 -128
rect -197 -130 -195 -128
rect -103 -130 -101 -128
rect -64 -130 -62 -128
rect 31 -130 33 -128
rect 41 -130 43 -128
rect 65 -130 67 -128
rect 76 -130 78 -128
rect 88 -130 90 -128
rect 182 -130 184 -128
rect 221 -130 223 -128
rect 316 -130 318 -128
rect 326 -130 328 -128
rect 350 -130 352 -128
rect 361 -130 363 -128
rect 373 -130 375 -128
rect 488 -130 490 -128
rect 657 -130 659 -128
rect 739 -141 741 -139
rect -688 -169 -686 -167
rect -673 -166 -671 -164
rect -663 -169 -661 -167
rect -647 -166 -645 -164
rect -634 -160 -632 -158
rect -617 -162 -615 -160
rect -626 -177 -624 -175
rect -593 -167 -591 -165
rect -580 -160 -578 -158
rect -563 -162 -561 -160
rect -572 -177 -570 -175
rect -539 -167 -537 -165
rect -529 -166 -527 -164
rect -505 -161 -503 -159
rect -513 -174 -511 -172
rect -494 -166 -492 -164
rect -470 -159 -468 -157
rect -482 -174 -480 -172
rect -454 -160 -452 -158
rect -437 -161 -435 -159
rect -446 -177 -444 -175
rect -413 -163 -411 -161
rect -403 -169 -401 -167
rect -388 -166 -386 -164
rect -378 -169 -376 -167
rect -362 -166 -360 -164
rect -349 -160 -347 -158
rect -332 -162 -330 -160
rect -341 -177 -339 -175
rect -308 -167 -306 -165
rect -295 -160 -293 -158
rect -278 -162 -276 -160
rect -287 -177 -285 -175
rect -254 -167 -252 -165
rect -244 -166 -242 -164
rect -220 -161 -218 -159
rect -228 -174 -226 -172
rect -209 -166 -207 -164
rect -185 -159 -183 -157
rect -197 -174 -195 -172
rect -169 -160 -167 -158
rect -152 -161 -150 -159
rect -161 -177 -159 -175
rect -128 -163 -126 -161
rect -118 -169 -116 -167
rect -103 -166 -101 -164
rect -93 -169 -91 -167
rect -77 -166 -75 -164
rect -64 -160 -62 -158
rect -47 -162 -45 -160
rect -56 -177 -54 -175
rect -23 -167 -21 -165
rect -10 -160 -8 -158
rect 7 -162 9 -160
rect -2 -177 0 -175
rect 31 -167 33 -165
rect 41 -166 43 -164
rect 65 -161 67 -159
rect 57 -174 59 -172
rect 76 -166 78 -164
rect 100 -159 102 -157
rect 88 -174 90 -172
rect 116 -160 118 -158
rect 133 -161 135 -159
rect 124 -177 126 -175
rect 157 -163 159 -161
rect 167 -169 169 -167
rect 182 -166 184 -164
rect 192 -169 194 -167
rect 208 -166 210 -164
rect 221 -160 223 -158
rect 238 -162 240 -160
rect 229 -177 231 -175
rect 262 -167 264 -165
rect 275 -160 277 -158
rect 292 -162 294 -160
rect 283 -177 285 -175
rect 316 -167 318 -165
rect 326 -166 328 -164
rect 350 -161 352 -159
rect 342 -174 344 -172
rect 361 -166 363 -164
rect 385 -159 387 -157
rect 373 -174 375 -172
rect 401 -160 403 -158
rect 418 -161 420 -159
rect 409 -177 411 -175
rect 442 -163 444 -161
rect 488 -161 490 -159
rect 470 -176 472 -174
rect 499 -177 501 -175
rect 460 -181 462 -179
rect 580 -161 582 -159
rect 535 -164 537 -162
rect 657 -152 659 -150
rect 705 -152 707 -150
rect 562 -176 564 -174
rect 591 -177 593 -175
rect 552 -182 554 -180
rect 705 -160 707 -158
rect 713 -160 715 -158
rect 713 -168 715 -166
rect 721 -168 723 -166
rect -733 -209 -731 -207
rect -688 -249 -686 -247
rect -673 -252 -671 -250
rect -663 -249 -661 -247
rect -626 -241 -624 -239
rect -647 -252 -645 -250
rect -634 -258 -632 -256
rect -617 -256 -615 -254
rect -572 -241 -570 -239
rect -593 -251 -591 -249
rect -580 -258 -578 -256
rect -563 -256 -561 -254
rect -513 -244 -511 -242
rect -539 -251 -537 -249
rect -529 -252 -527 -250
rect -482 -244 -480 -242
rect -494 -252 -492 -250
rect -505 -257 -503 -255
rect -446 -241 -444 -239
rect -470 -259 -468 -257
rect -454 -258 -452 -256
rect -403 -249 -401 -247
rect -413 -255 -411 -253
rect -437 -257 -435 -255
rect -388 -252 -386 -250
rect -378 -249 -376 -247
rect -341 -241 -339 -239
rect -362 -252 -360 -250
rect -349 -258 -347 -256
rect -332 -256 -330 -254
rect -287 -241 -285 -239
rect -308 -251 -306 -249
rect -295 -258 -293 -256
rect -278 -256 -276 -254
rect -228 -244 -226 -242
rect -254 -251 -252 -249
rect -244 -252 -242 -250
rect -197 -244 -195 -242
rect -209 -252 -207 -250
rect -220 -257 -218 -255
rect -161 -241 -159 -239
rect -185 -259 -183 -257
rect -169 -258 -167 -256
rect -118 -249 -116 -247
rect -128 -255 -126 -253
rect -152 -257 -150 -255
rect -103 -252 -101 -250
rect -93 -249 -91 -247
rect -56 -241 -54 -239
rect -77 -252 -75 -250
rect -64 -258 -62 -256
rect -47 -256 -45 -254
rect -2 -241 0 -239
rect -23 -251 -21 -249
rect -10 -258 -8 -256
rect 7 -256 9 -254
rect 57 -244 59 -242
rect 31 -251 33 -249
rect 41 -252 43 -250
rect 88 -244 90 -242
rect 76 -252 78 -250
rect 65 -257 67 -255
rect 124 -241 126 -239
rect 100 -259 102 -257
rect 116 -258 118 -256
rect 167 -249 169 -247
rect 157 -255 159 -253
rect 133 -257 135 -255
rect 182 -252 184 -250
rect 192 -249 194 -247
rect 229 -241 231 -239
rect 208 -252 210 -250
rect 221 -258 223 -256
rect 238 -256 240 -254
rect 283 -241 285 -239
rect 262 -251 264 -249
rect 275 -258 277 -256
rect 292 -256 294 -254
rect 342 -244 344 -242
rect 316 -251 318 -249
rect 326 -252 328 -250
rect 373 -244 375 -242
rect 361 -252 363 -250
rect 350 -257 352 -255
rect 409 -241 411 -239
rect 385 -259 387 -257
rect 401 -258 403 -256
rect 460 -237 462 -235
rect 470 -242 472 -240
rect 493 -241 495 -239
rect 442 -255 444 -253
rect 418 -257 420 -255
rect 482 -257 484 -255
rect 554 -237 556 -235
rect 562 -243 564 -241
rect 599 -241 601 -239
rect 572 -257 574 -255
rect 739 -277 741 -275
rect -673 -288 -671 -286
rect -634 -288 -632 -286
rect -539 -288 -537 -286
rect -529 -288 -527 -286
rect -505 -288 -503 -286
rect -494 -288 -492 -286
rect -482 -288 -480 -286
rect -388 -288 -386 -286
rect -349 -288 -347 -286
rect -254 -288 -252 -286
rect -244 -288 -242 -286
rect -220 -288 -218 -286
rect -209 -288 -207 -286
rect -197 -288 -195 -286
rect -103 -288 -101 -286
rect -64 -288 -62 -286
rect 31 -288 33 -286
rect 41 -288 43 -286
rect 65 -288 67 -286
rect 76 -288 78 -286
rect 88 -288 90 -286
rect 182 -288 184 -286
rect 221 -288 223 -286
rect 316 -288 318 -286
rect 326 -288 328 -286
rect 350 -288 352 -286
rect 361 -288 363 -286
rect 373 -288 375 -286
rect 460 -289 462 -287
rect 681 -289 683 -287
rect -688 -296 -686 -294
rect -580 -296 -578 -294
rect -513 -296 -511 -294
rect -470 -296 -468 -294
rect -454 -296 -452 -294
rect -403 -296 -401 -294
rect -295 -296 -293 -294
rect -228 -296 -226 -294
rect -185 -296 -183 -294
rect -169 -296 -167 -294
rect -118 -296 -116 -294
rect -10 -296 -8 -294
rect 57 -296 59 -294
rect 100 -296 102 -294
rect 116 -296 118 -294
rect 167 -296 169 -294
rect 275 -296 277 -294
rect 342 -296 344 -294
rect 385 -296 387 -294
rect 401 -296 403 -294
rect 442 -297 444 -295
rect 554 -297 556 -295
rect 562 -297 564 -295
rect 657 -297 659 -295
rect -698 -304 -696 -302
rect -663 -304 -661 -302
rect -647 -304 -645 -302
rect -626 -304 -624 -302
rect -572 -304 -570 -302
rect -362 -304 -360 -302
rect -341 -304 -339 -302
rect -287 -304 -285 -302
rect -77 -304 -75 -302
rect -56 -304 -54 -302
rect -2 -304 0 -302
rect 208 -304 210 -302
rect 229 -304 231 -302
rect 283 -304 285 -302
rect 470 -305 472 -303
rect 689 -305 691 -303
rect -593 -312 -591 -310
rect -482 -312 -480 -310
rect -308 -312 -306 -310
rect -197 -312 -195 -310
rect -23 -312 -21 -310
rect 88 -312 90 -310
rect 262 -312 264 -310
rect 373 -312 375 -310
rect 482 -313 484 -311
rect 697 -313 699 -311
rect -663 -320 -661 -318
rect -446 -320 -444 -318
rect -378 -320 -376 -318
rect -161 -320 -159 -318
rect -93 -320 -91 -318
rect 124 -320 126 -318
rect 192 -320 194 -318
rect 409 -320 411 -318
rect 572 -321 574 -319
rect 705 -321 707 -319
rect -617 -328 -615 -326
rect -563 -328 -561 -326
rect -437 -328 -435 -326
rect -332 -328 -330 -326
rect -278 -328 -276 -326
rect -152 -328 -150 -326
rect -47 -328 -45 -326
rect 7 -328 9 -326
rect 133 -328 135 -326
rect 157 -328 159 -326
rect 200 -328 202 -326
rect 238 -328 240 -326
rect 292 -328 294 -326
rect 418 -328 420 -326
rect 599 -329 601 -327
rect 713 -329 715 -327
rect -617 -336 -615 -334
rect -332 -336 -330 -334
rect -47 -336 -45 -334
rect 238 -336 240 -334
rect 633 -337 635 -335
rect -663 -344 -661 -342
rect -378 -344 -376 -342
rect -93 -344 -91 -342
rect 192 -344 194 -342
rect 200 -344 202 -342
rect 493 -344 495 -342
rect -706 -352 -704 -350
rect -403 -352 -401 -350
rect -128 -352 -126 -350
rect 158 -352 160 -350
rect 167 -352 169 -350
rect 641 -352 643 -350
rect -714 -360 -712 -358
rect -688 -360 -686 -358
rect -118 -360 -116 -358
rect 649 -360 651 -358
rect -413 -369 -411 -367
rect 665 -369 667 -367
rect 158 -377 160 -375
rect 673 -377 675 -375
<< labels >>
rlabel alu1 540 138 540 138 6 vdd
rlabel alu1 480 138 480 138 6 vdd
rlabel alu1 590 138 590 138 6 vdd
rlabel via1 561 63 561 63 1 En
rlabel alu1 540 146 540 146 8 vdd
rlabel alu1 480 146 480 146 8 vdd
rlabel alu1 590 146 590 146 8 vdd
rlabel via1 598 229 598 229 1 A1
rlabel via1 598 55 598 55 1 A0
rlabel via1 456 253 456 253 5 Y2
rlabel via1 516 253 516 253 5 Y0
rlabel via1 516 47 516 47 1 Y3
rlabel via1 456 47 456 47 1 Y1
rlabel alu1 573 210 573 210 1 vss
rlabel alu1 508 210 508 210 1 vss
rlabel alu1 462 210 462 210 1 vss
rlabel alu1 573 74 573 74 1 vss
rlabel alu1 523 74 523 74 1 vss
rlabel alu1 463 74 463 74 1 vss
rlabel alu1 588 -204 588 -204 2 vdd
rlabel alu1 588 -140 588 -140 2 vss
rlabel alu1 496 -204 496 -204 2 vdd
rlabel alu1 496 -140 496 -140 2 vss
rlabel alu1 588 -212 588 -212 4 vdd
rlabel alu1 588 -276 588 -276 4 vss
rlabel alu1 496 -212 496 -212 4 vdd
rlabel alu1 496 -276 496 -276 4 vss
rlabel via1 -697 -303 -697 -303 1 RorW
rlabel via1 -705 -351 -705 -351 1 In2
rlabel via1 642 -351 642 -351 1 In0
rlabel via1 650 -359 650 -359 1 In1
rlabel via1 -713 -359 -713 -359 1 In3
rlabel via1 536 -163 536 -163 1 D3
rlabel alu1 628 -163 628 -163 1 D2
rlabel alu1 536 -246 536 -246 1 D1
rlabel alu1 628 -245 628 -245 1 D0
rlabel via1 561 221 561 221 1 En
<< end >>
