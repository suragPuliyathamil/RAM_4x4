magic
tech scmos
timestamp 1607485093
<< ab >>
rect -13 -5 19 67
rect 22 -5 54 67
<< nwell >>
rect -18 27 59 72
<< pwell >>
rect -18 -10 59 27
<< poly >>
rect -2 61 0 65
rect 5 61 7 65
rect 33 61 35 65
rect 40 61 42 65
rect -2 27 0 33
rect 5 30 7 33
rect -6 25 0 27
rect -6 23 -4 25
rect -2 23 0 25
rect 4 28 10 30
rect 4 26 6 28
rect 8 26 10 28
rect 33 27 35 33
rect 40 30 42 33
rect 4 24 10 26
rect 29 25 35 27
rect -6 21 0 23
rect -4 18 -2 21
rect 7 15 9 24
rect 29 23 31 25
rect 33 23 35 25
rect 39 28 45 30
rect 39 26 41 28
rect 43 26 45 28
rect 39 24 45 26
rect 29 21 35 23
rect 31 18 33 21
rect -4 6 -2 10
rect 42 15 44 24
rect 7 2 9 7
rect 31 6 33 10
rect 42 2 44 7
<< ndif >>
rect -11 14 -4 18
rect -11 12 -9 14
rect -7 12 -4 14
rect -11 10 -4 12
rect -2 15 3 18
rect -2 11 7 15
rect -2 10 2 11
rect 0 9 2 10
rect 4 9 7 11
rect 0 7 7 9
rect 9 7 17 15
rect 24 14 31 18
rect 24 12 26 14
rect 28 12 31 14
rect 24 10 31 12
rect 33 15 38 18
rect 33 11 42 15
rect 33 10 37 11
rect 11 2 17 7
rect 35 9 37 10
rect 39 9 42 11
rect 35 7 42 9
rect 44 7 52 15
rect 11 0 13 2
rect 15 0 17 2
rect 11 -2 17 0
rect 46 2 52 7
rect 46 0 48 2
rect 50 0 52 2
rect 46 -2 52 0
<< pdif >>
rect -11 59 -2 61
rect -11 57 -9 59
rect -7 57 -2 59
rect -11 52 -2 57
rect -11 50 -9 52
rect -7 50 -2 52
rect -11 33 -2 50
rect 0 33 5 61
rect 7 54 12 61
rect 24 59 33 61
rect 24 57 26 59
rect 28 57 33 59
rect 7 52 14 54
rect 7 50 10 52
rect 12 50 14 52
rect 7 45 14 50
rect 7 43 10 45
rect 12 43 14 45
rect 7 41 14 43
rect 24 52 33 57
rect 24 50 26 52
rect 28 50 33 52
rect 7 33 12 41
rect 24 33 33 50
rect 35 33 40 61
rect 42 54 47 61
rect 42 52 49 54
rect 42 50 45 52
rect 47 50 49 52
rect 42 45 49 50
rect 42 43 45 45
rect 47 43 49 45
rect 42 41 49 43
rect 42 33 47 41
<< alu1 >>
rect -15 59 56 67
rect 8 52 14 53
rect 8 50 10 52
rect 12 50 14 52
rect 8 46 14 50
rect 43 52 49 53
rect 43 50 45 52
rect 47 50 49 52
rect 43 46 49 50
rect 8 45 17 46
rect 8 43 10 45
rect 12 43 17 45
rect 8 42 17 43
rect 43 45 52 46
rect 43 43 45 45
rect 47 43 52 45
rect 43 42 52 43
rect -3 34 1 38
rect -3 33 9 34
rect -3 31 6 33
rect 8 31 9 33
rect -3 30 9 31
rect -11 26 -7 30
rect 5 28 9 30
rect 5 26 6 28
rect 8 26 9 28
rect -11 25 1 26
rect -11 23 -10 25
rect -8 23 -4 25
rect -2 23 1 25
rect 5 24 9 26
rect -11 22 1 23
rect -3 16 1 22
rect 13 20 17 42
rect 32 34 36 38
rect 32 33 44 34
rect 32 31 37 33
rect 39 31 44 33
rect 32 30 44 31
rect 24 26 28 30
rect 40 28 44 30
rect 40 26 41 28
rect 43 26 44 28
rect 24 25 36 26
rect 24 23 25 25
rect 27 23 31 25
rect 33 23 36 25
rect 40 24 44 26
rect 24 22 36 23
rect 13 18 14 20
rect 16 18 17 20
rect 13 14 17 18
rect 32 16 36 22
rect 48 18 52 42
rect 48 16 49 18
rect 51 16 52 18
rect 5 12 17 14
rect 0 11 17 12
rect 0 9 2 11
rect 4 9 17 11
rect 0 8 17 9
rect 48 14 52 16
rect 40 12 52 14
rect 35 11 52 12
rect 35 9 37 11
rect 39 9 52 11
rect 35 8 52 9
rect -15 2 56 3
rect -15 0 -8 2
rect -6 0 13 2
rect 15 0 27 2
rect 29 0 48 2
rect 50 0 56 2
rect -15 -5 56 0
rect -11 -11 -7 -10
rect -11 -13 -10 -11
rect -8 -13 -7 -11
rect -11 -14 -7 -13
rect 13 -11 28 -10
rect 13 -13 14 -11
rect 16 -13 25 -11
rect 27 -13 28 -11
rect 13 -14 28 -13
rect 36 -11 40 -10
rect 36 -13 37 -11
rect 39 -13 40 -11
rect 36 -14 40 -13
rect 5 -19 52 -18
rect 5 -21 6 -19
rect 8 -21 49 -19
rect 51 -21 52 -19
rect 5 -22 52 -21
<< alu2 >>
rect 5 33 9 34
rect 5 31 6 33
rect 8 31 9 33
rect -11 25 -7 26
rect -11 23 -10 25
rect -8 23 -7 25
rect -11 -11 -7 23
rect -11 -13 -10 -11
rect -8 -13 -7 -11
rect -11 -14 -7 -13
rect 5 -19 9 31
rect 36 33 40 34
rect 36 31 37 33
rect 39 31 40 33
rect 24 25 28 26
rect 24 23 25 25
rect 27 23 28 25
rect 13 20 17 21
rect 13 18 14 20
rect 16 18 17 20
rect 13 -11 17 18
rect 13 -13 14 -11
rect 16 -13 17 -11
rect 13 -14 17 -13
rect 24 -11 28 23
rect 24 -13 25 -11
rect 27 -13 28 -11
rect 24 -14 28 -13
rect 36 -11 40 31
rect 36 -13 37 -11
rect 39 -13 40 -11
rect 36 -14 40 -13
rect 48 18 52 19
rect 48 16 49 18
rect 51 16 52 18
rect 5 -21 6 -19
rect 8 -21 9 -19
rect 5 -22 9 -21
rect 48 -19 52 16
rect 48 -21 49 -19
rect 51 -21 52 -19
rect 48 -22 52 -21
<< ptie >>
rect -10 2 -4 4
rect -10 0 -8 2
rect -6 0 -4 2
rect -10 -2 -4 0
rect 25 2 31 4
rect 25 0 27 2
rect 29 0 31 2
rect 25 -2 31 0
<< nmos >>
rect -4 10 -2 18
rect 7 7 9 15
rect 31 10 33 18
rect 42 7 44 15
<< pmos >>
rect -2 33 0 61
rect 5 33 7 61
rect 33 33 35 61
rect 40 33 42 61
<< polyct1 >>
rect -4 23 -2 25
rect 6 26 8 28
rect 31 23 33 25
rect 41 26 43 28
<< ndifct0 >>
rect -9 12 -7 14
rect 26 12 28 14
<< ndifct1 >>
rect 2 9 4 11
rect 37 9 39 11
rect 13 0 15 2
rect 48 0 50 2
<< ptiect1 >>
rect -8 0 -6 2
rect 27 0 29 2
<< pdifct0 >>
rect -9 57 -7 59
rect -9 50 -7 52
rect 26 57 28 59
rect 26 50 28 52
<< pdifct1 >>
rect 10 50 12 52
rect 10 43 12 45
rect 45 50 47 52
rect 45 43 47 45
<< alu0 >>
rect -10 57 -9 59
rect -7 57 -6 59
rect -10 52 -6 57
rect 25 57 26 59
rect 28 57 29 59
rect -10 50 -9 52
rect -7 50 -6 52
rect -10 48 -6 50
rect 25 52 29 57
rect 25 50 26 52
rect 28 50 29 52
rect 25 48 29 50
rect -10 14 -6 16
rect -10 12 -9 14
rect -7 12 -6 14
rect -10 3 -6 12
rect 25 14 29 16
rect 25 12 26 14
rect 28 12 29 14
rect 25 3 29 12
<< via1 >>
rect 6 31 8 33
rect -10 23 -8 25
rect 37 31 39 33
rect 25 23 27 25
rect 14 18 16 20
rect 49 16 51 18
rect -10 -13 -8 -11
rect 14 -13 16 -11
rect 25 -13 27 -11
rect 37 -13 39 -11
rect 6 -21 8 -19
rect 49 -21 51 -19
<< labels >>
rlabel alu1 3 -1 3 -1 4 vss
rlabel alu1 3 63 3 63 4 vdd
rlabel alu1 38 63 38 63 4 vdd
rlabel alu1 38 -1 38 -1 4 vss
rlabel via1 15 -12 15 -12 1 Q_bar
rlabel via1 50 -20 50 -20 1 Q
rlabel via1 -9 -12 -9 -12 1 S
rlabel via1 38 -12 38 -12 1 R
<< end >>
