magic
tech scmos
timestamp 1607528933
<< ab >>
rect -133 -117 -109 27
rect -99 -73 -43 27
rect -99 -109 -75 -73
rect -74 -109 -43 -73
rect -99 -117 -43 -109
rect -39 19 17 27
rect -39 -17 -15 19
rect -14 -17 17 19
rect -39 -73 17 -17
rect -39 -117 -15 -73
rect -14 -117 17 -73
<< nwell >>
rect -138 -85 22 -5
<< pwell >>
rect -138 -5 22 32
rect -138 -122 22 -85
<< poly >>
rect -81 15 -79 20
rect -74 15 -72 20
rect -67 15 -65 20
rect -120 10 -118 15
rect -54 11 -52 16
rect -21 15 -19 20
rect -14 15 -12 20
rect -7 15 -5 20
rect 6 11 8 16
rect -120 -2 -118 1
rect -81 -2 -79 2
rect -124 -4 -118 -2
rect -124 -6 -122 -4
rect -120 -6 -118 -4
rect -124 -8 -118 -6
rect -90 -4 -79 -2
rect -90 -6 -88 -4
rect -86 -6 -84 -4
rect -90 -8 -84 -6
rect -120 -11 -118 -8
rect -86 -17 -84 -8
rect -74 -9 -72 2
rect -67 -2 -65 2
rect -54 -2 -52 2
rect -21 -2 -19 2
rect -68 -4 -62 -2
rect -68 -6 -66 -4
rect -64 -6 -62 -4
rect -68 -8 -62 -6
rect -58 -4 -52 -2
rect -58 -6 -56 -4
rect -54 -6 -52 -4
rect -58 -8 -52 -6
rect -30 -4 -19 -2
rect -30 -6 -28 -4
rect -26 -6 -24 -4
rect -30 -8 -24 -6
rect -78 -11 -72 -9
rect -78 -13 -76 -11
rect -74 -13 -72 -11
rect -78 -15 -72 -13
rect -120 -34 -118 -29
rect -74 -18 -72 -15
rect -64 -18 -62 -8
rect -54 -13 -52 -8
rect -86 -35 -84 -30
rect -26 -17 -24 -8
rect -14 -9 -12 2
rect -7 -2 -5 2
rect 6 -2 8 2
rect -8 -4 -2 -2
rect -8 -6 -6 -4
rect -4 -6 -2 -4
rect -8 -8 -2 -6
rect 2 -4 8 -2
rect 2 -6 4 -4
rect 6 -6 8 -4
rect 2 -8 8 -6
rect -18 -11 -12 -9
rect -18 -13 -16 -11
rect -14 -13 -12 -11
rect -18 -15 -12 -13
rect -14 -18 -12 -15
rect -4 -18 -2 -8
rect 6 -13 8 -8
rect -74 -36 -72 -31
rect -64 -36 -62 -31
rect -54 -36 -52 -31
rect -26 -35 -24 -30
rect -14 -36 -12 -31
rect -4 -36 -2 -31
rect 6 -36 8 -31
rect -120 -61 -118 -56
rect -86 -60 -84 -55
rect -74 -59 -72 -54
rect -64 -59 -62 -54
rect -54 -59 -52 -54
rect -120 -82 -118 -79
rect -86 -82 -84 -73
rect -74 -75 -72 -72
rect -78 -77 -72 -75
rect -78 -79 -76 -77
rect -74 -79 -72 -77
rect -78 -81 -72 -79
rect -124 -84 -118 -82
rect -124 -86 -122 -84
rect -120 -86 -118 -84
rect -124 -88 -118 -86
rect -90 -84 -84 -82
rect -90 -86 -88 -84
rect -86 -86 -84 -84
rect -90 -88 -79 -86
rect -120 -91 -118 -88
rect -81 -92 -79 -88
rect -74 -92 -72 -81
rect -64 -82 -62 -72
rect -26 -60 -24 -55
rect -14 -59 -12 -54
rect -4 -59 -2 -54
rect 6 -59 8 -54
rect -54 -82 -52 -77
rect -26 -82 -24 -73
rect -14 -75 -12 -72
rect -18 -77 -12 -75
rect -18 -79 -16 -77
rect -14 -79 -12 -77
rect -18 -81 -12 -79
rect -68 -84 -62 -82
rect -68 -86 -66 -84
rect -64 -86 -62 -84
rect -68 -88 -62 -86
rect -58 -84 -52 -82
rect -58 -86 -56 -84
rect -54 -86 -52 -84
rect -58 -88 -52 -86
rect -30 -84 -24 -82
rect -30 -86 -28 -84
rect -26 -86 -24 -84
rect -30 -88 -19 -86
rect -67 -92 -65 -88
rect -54 -92 -52 -88
rect -21 -92 -19 -88
rect -14 -92 -12 -81
rect -4 -82 -2 -72
rect 6 -82 8 -77
rect -8 -84 -2 -82
rect -8 -86 -6 -84
rect -4 -86 -2 -84
rect -8 -88 -2 -86
rect 2 -84 8 -82
rect 2 -86 4 -84
rect 6 -86 8 -84
rect 2 -88 8 -86
rect -7 -92 -5 -88
rect 6 -92 8 -88
rect -120 -105 -118 -100
rect -81 -110 -79 -105
rect -74 -110 -72 -105
rect -67 -110 -65 -105
rect -54 -106 -52 -101
rect -21 -110 -19 -105
rect -14 -110 -12 -105
rect -7 -110 -5 -105
rect 6 -106 8 -101
<< ndif >>
rect -63 22 -56 24
rect -63 20 -60 22
rect -58 20 -56 22
rect -63 15 -56 20
rect -3 22 4 24
rect -3 20 0 22
rect 2 20 4 22
rect -88 13 -81 15
rect -88 11 -86 13
rect -84 11 -81 13
rect -131 8 -120 10
rect -131 6 -129 8
rect -127 6 -120 8
rect -131 1 -120 6
rect -118 7 -113 10
rect -88 9 -81 11
rect -118 5 -111 7
rect -118 3 -115 5
rect -113 3 -111 5
rect -118 1 -111 3
rect -86 2 -81 9
rect -79 2 -74 15
rect -72 2 -67 15
rect -65 11 -56 15
rect -3 15 4 20
rect -28 13 -21 15
rect -28 11 -26 13
rect -24 11 -21 13
rect -65 2 -54 11
rect -52 8 -47 11
rect -28 9 -21 11
rect -52 6 -45 8
rect -52 4 -49 6
rect -47 4 -45 6
rect -52 2 -45 4
rect -26 2 -21 9
rect -19 2 -14 15
rect -12 2 -7 15
rect -5 11 4 15
rect -5 2 6 11
rect 8 8 13 11
rect 8 6 15 8
rect 8 4 11 6
rect 13 4 15 6
rect 8 2 15 4
rect -131 -96 -120 -91
rect -131 -98 -129 -96
rect -127 -98 -120 -96
rect -131 -100 -120 -98
rect -118 -93 -111 -91
rect -118 -95 -115 -93
rect -113 -95 -111 -93
rect -118 -97 -111 -95
rect -118 -100 -113 -97
rect -86 -99 -81 -92
rect -88 -101 -81 -99
rect -88 -103 -86 -101
rect -84 -103 -81 -101
rect -88 -105 -81 -103
rect -79 -105 -74 -92
rect -72 -105 -67 -92
rect -65 -101 -54 -92
rect -52 -94 -45 -92
rect -52 -96 -49 -94
rect -47 -96 -45 -94
rect -52 -98 -45 -96
rect -52 -101 -47 -98
rect -26 -99 -21 -92
rect -28 -101 -21 -99
rect -65 -105 -56 -101
rect -63 -110 -56 -105
rect -28 -103 -26 -101
rect -24 -103 -21 -101
rect -28 -105 -21 -103
rect -19 -105 -14 -92
rect -12 -105 -7 -92
rect -5 -101 6 -92
rect 8 -94 15 -92
rect 8 -96 11 -94
rect 13 -96 15 -94
rect 8 -98 15 -96
rect 8 -101 13 -98
rect -5 -105 4 -101
rect -63 -112 -60 -110
rect -58 -112 -56 -110
rect -63 -114 -56 -112
rect -3 -110 4 -105
rect -3 -112 0 -110
rect 2 -112 4 -110
rect -3 -114 4 -112
<< pdif >>
rect -129 -28 -120 -11
rect -129 -30 -126 -28
rect -124 -29 -120 -28
rect -118 -13 -111 -11
rect -118 -15 -115 -13
rect -113 -15 -111 -13
rect -118 -20 -111 -15
rect -118 -22 -115 -20
rect -113 -22 -111 -20
rect -118 -24 -111 -22
rect -93 -19 -86 -17
rect -93 -21 -91 -19
rect -89 -21 -86 -19
rect -118 -29 -113 -24
rect -93 -26 -86 -21
rect -93 -28 -91 -26
rect -89 -28 -86 -26
rect -124 -30 -122 -29
rect -129 -32 -122 -30
rect -93 -30 -86 -28
rect -84 -18 -79 -17
rect -60 -18 -54 -13
rect -84 -30 -74 -18
rect -82 -31 -74 -30
rect -72 -20 -64 -18
rect -72 -22 -69 -20
rect -67 -22 -64 -20
rect -72 -27 -64 -22
rect -72 -29 -69 -27
rect -67 -29 -64 -27
rect -72 -31 -64 -29
rect -62 -27 -54 -18
rect -62 -29 -59 -27
rect -57 -29 -54 -27
rect -62 -31 -54 -29
rect -52 -15 -45 -13
rect -52 -17 -49 -15
rect -47 -17 -45 -15
rect -52 -22 -45 -17
rect -52 -24 -49 -22
rect -47 -24 -45 -22
rect -52 -26 -45 -24
rect -33 -19 -26 -17
rect -33 -21 -31 -19
rect -29 -21 -26 -19
rect -33 -26 -26 -21
rect -52 -31 -47 -26
rect -33 -28 -31 -26
rect -29 -28 -26 -26
rect -33 -30 -26 -28
rect -24 -18 -19 -17
rect 0 -18 6 -13
rect -24 -30 -14 -18
rect -82 -38 -76 -31
rect -22 -31 -14 -30
rect -12 -20 -4 -18
rect -12 -22 -9 -20
rect -7 -22 -4 -20
rect -12 -27 -4 -22
rect -12 -29 -9 -27
rect -7 -29 -4 -27
rect -12 -31 -4 -29
rect -2 -27 6 -18
rect -2 -29 1 -27
rect 3 -29 6 -27
rect -2 -31 6 -29
rect 8 -15 15 -13
rect 8 -17 11 -15
rect 13 -17 15 -15
rect 8 -22 15 -17
rect 8 -24 11 -22
rect 13 -24 15 -22
rect 8 -26 15 -24
rect 8 -31 13 -26
rect -82 -40 -80 -38
rect -78 -40 -76 -38
rect -82 -42 -76 -40
rect -22 -38 -16 -31
rect -22 -40 -20 -38
rect -18 -40 -16 -38
rect -22 -42 -16 -40
rect -82 -50 -76 -48
rect -82 -52 -80 -50
rect -78 -52 -76 -50
rect -129 -60 -122 -58
rect -129 -62 -126 -60
rect -124 -61 -122 -60
rect -82 -59 -76 -52
rect -22 -50 -16 -48
rect -22 -52 -20 -50
rect -18 -52 -16 -50
rect -82 -60 -74 -59
rect -124 -62 -120 -61
rect -129 -79 -120 -62
rect -118 -66 -113 -61
rect -93 -62 -86 -60
rect -93 -64 -91 -62
rect -89 -64 -86 -62
rect -118 -68 -111 -66
rect -118 -70 -115 -68
rect -113 -70 -111 -68
rect -118 -75 -111 -70
rect -93 -69 -86 -64
rect -93 -71 -91 -69
rect -89 -71 -86 -69
rect -93 -73 -86 -71
rect -84 -72 -74 -60
rect -72 -61 -64 -59
rect -72 -63 -69 -61
rect -67 -63 -64 -61
rect -72 -68 -64 -63
rect -72 -70 -69 -68
rect -67 -70 -64 -68
rect -72 -72 -64 -70
rect -62 -61 -54 -59
rect -62 -63 -59 -61
rect -57 -63 -54 -61
rect -62 -72 -54 -63
rect -84 -73 -79 -72
rect -118 -77 -115 -75
rect -113 -77 -111 -75
rect -118 -79 -111 -77
rect -60 -77 -54 -72
rect -52 -64 -47 -59
rect -22 -59 -16 -52
rect -22 -60 -14 -59
rect -33 -62 -26 -60
rect -33 -64 -31 -62
rect -29 -64 -26 -62
rect -52 -66 -45 -64
rect -52 -68 -49 -66
rect -47 -68 -45 -66
rect -52 -73 -45 -68
rect -33 -69 -26 -64
rect -33 -71 -31 -69
rect -29 -71 -26 -69
rect -33 -73 -26 -71
rect -24 -72 -14 -60
rect -12 -61 -4 -59
rect -12 -63 -9 -61
rect -7 -63 -4 -61
rect -12 -68 -4 -63
rect -12 -70 -9 -68
rect -7 -70 -4 -68
rect -12 -72 -4 -70
rect -2 -61 6 -59
rect -2 -63 1 -61
rect 3 -63 6 -61
rect -2 -72 6 -63
rect -24 -73 -19 -72
rect -52 -75 -49 -73
rect -47 -75 -45 -73
rect -52 -77 -45 -75
rect 0 -77 6 -72
rect 8 -64 13 -59
rect 8 -66 15 -64
rect 8 -68 11 -66
rect 13 -68 15 -66
rect 8 -73 15 -68
rect 8 -75 11 -73
rect 13 -75 15 -73
rect 8 -77 15 -75
<< alu1 >>
rect -49 67 -45 68
rect -49 65 -48 67
rect -46 65 -45 67
rect -49 64 -45 65
rect 11 67 15 68
rect 11 65 12 67
rect 14 65 15 67
rect 11 64 15 65
rect -143 59 -9 60
rect -143 57 -142 59
rect -140 57 -72 59
rect -70 57 -12 59
rect -10 57 -9 59
rect -143 56 -9 57
rect -159 51 -81 52
rect -159 49 -158 51
rect -156 49 -114 51
rect -112 49 -84 51
rect -82 49 -81 51
rect -159 48 -81 49
rect -151 43 -19 44
rect -151 41 -150 43
rect -148 41 -130 43
rect -128 41 -22 43
rect -20 41 -19 43
rect -151 40 -19 41
rect -94 35 -30 36
rect -94 33 -93 35
rect -91 33 -33 35
rect -31 33 -30 35
rect -94 32 -30 33
rect -135 24 29 27
rect -135 22 25 24
rect 27 22 29 24
rect -135 20 -128 22
rect -126 20 -116 22
rect -114 20 -60 22
rect -58 20 -50 22
rect -48 20 0 22
rect 2 20 10 22
rect 12 20 29 22
rect -135 19 29 20
rect -115 12 -111 14
rect -115 10 -114 12
rect -112 10 -111 12
rect -123 -2 -119 6
rect -115 5 -111 10
rect -113 3 -111 5
rect -131 -4 -119 -2
rect -131 -6 -130 -4
rect -128 -6 -122 -4
rect -120 -6 -119 -4
rect -131 -8 -119 -6
rect -115 -13 -111 3
rect -90 5 -77 6
rect -90 3 -84 5
rect -82 3 -77 5
rect -90 0 -77 3
rect -73 5 -69 6
rect -73 3 -72 5
rect -70 3 -69 5
rect -90 -4 -84 0
rect -90 -6 -88 -4
rect -86 -6 -84 -4
rect -90 -7 -84 -6
rect -73 -3 -69 3
rect -49 6 -45 14
rect -47 4 -45 6
rect -73 -4 -60 -3
rect -73 -6 -66 -4
rect -64 -6 -60 -4
rect -73 -7 -60 -6
rect -113 -15 -111 -13
rect -94 -12 -76 -11
rect -94 -14 -93 -12
rect -91 -13 -76 -12
rect -74 -13 -68 -11
rect -91 -14 -68 -13
rect -94 -15 -68 -14
rect -49 0 -45 4
rect -31 3 -17 6
rect -31 1 -30 3
rect -28 1 -17 3
rect -31 0 -17 1
rect -13 5 -9 6
rect -13 3 -12 5
rect -10 3 -9 5
rect -49 -2 -48 0
rect -46 -2 -45 0
rect -115 -18 -111 -15
rect -123 -20 -111 -18
rect -123 -22 -115 -20
rect -113 -22 -111 -20
rect -123 -24 -111 -22
rect -82 -23 -76 -15
rect -49 -15 -45 -2
rect -30 -4 -24 0
rect -30 -6 -28 -4
rect -26 -6 -24 -4
rect -30 -7 -24 -6
rect -13 -3 -9 3
rect 11 6 15 14
rect 13 4 15 6
rect -13 -4 0 -3
rect -13 -6 -6 -4
rect -4 -6 0 -4
rect -13 -7 0 -6
rect -30 -12 -16 -11
rect -30 -14 -22 -12
rect -20 -13 -16 -12
rect -14 -13 -8 -11
rect -20 -14 -8 -13
rect -30 -15 -8 -14
rect 11 0 15 4
rect 11 -2 12 0
rect 14 -2 15 0
rect -47 -17 -45 -15
rect -49 -19 -45 -17
rect -58 -22 -45 -19
rect -58 -23 -49 -22
rect -50 -24 -49 -23
rect -47 -24 -45 -22
rect -50 -32 -45 -24
rect -22 -23 -16 -15
rect 11 -15 15 -2
rect 13 -17 15 -15
rect 11 -19 15 -17
rect 2 -22 15 -19
rect 2 -23 11 -22
rect 10 -24 11 -23
rect 13 -24 15 -22
rect 10 -32 15 -24
rect -135 -38 19 -37
rect -135 -40 -128 -38
rect -126 -40 -116 -38
rect -114 -40 -94 -38
rect -92 -40 -80 -38
rect -78 -40 -34 -38
rect -32 -40 -20 -38
rect -18 -40 19 -38
rect -135 -50 19 -40
rect -135 -52 -128 -50
rect -126 -52 -116 -50
rect -114 -52 -94 -50
rect -92 -52 -80 -50
rect -78 -52 -34 -50
rect -32 -52 -20 -50
rect -18 -52 19 -50
rect -135 -53 19 -52
rect -123 -68 -111 -66
rect -123 -70 -115 -68
rect -113 -70 -111 -68
rect -123 -72 -111 -70
rect -115 -75 -111 -72
rect -82 -75 -76 -67
rect -50 -66 -45 -58
rect -50 -67 -49 -66
rect -58 -68 -49 -67
rect -47 -68 -45 -66
rect -58 -71 -45 -68
rect -113 -77 -111 -75
rect -131 -84 -119 -82
rect -131 -86 -130 -84
rect -128 -86 -122 -84
rect -120 -86 -119 -84
rect -131 -88 -119 -86
rect -123 -96 -119 -88
rect -115 -93 -111 -77
rect -90 -76 -68 -75
rect -90 -78 -82 -76
rect -80 -77 -68 -76
rect -80 -78 -76 -77
rect -90 -79 -76 -78
rect -74 -79 -68 -77
rect -49 -73 -45 -71
rect -47 -75 -45 -73
rect -22 -75 -16 -67
rect 10 -66 15 -58
rect 10 -67 11 -66
rect 2 -68 11 -67
rect 13 -68 15 -66
rect 2 -71 15 -68
rect -90 -84 -84 -83
rect -90 -86 -88 -84
rect -86 -86 -84 -84
rect -90 -90 -84 -86
rect -73 -84 -60 -83
rect -73 -86 -66 -84
rect -64 -86 -60 -84
rect -73 -87 -60 -86
rect -113 -95 -111 -93
rect -115 -100 -111 -95
rect -91 -91 -77 -90
rect -91 -93 -90 -91
rect -88 -93 -77 -91
rect -91 -96 -77 -93
rect -73 -93 -69 -87
rect -49 -86 -45 -75
rect -30 -76 -8 -75
rect -30 -78 -22 -76
rect -20 -77 -8 -76
rect -20 -78 -16 -77
rect -30 -79 -16 -78
rect -14 -79 -8 -77
rect 11 -73 15 -71
rect 13 -75 15 -73
rect -49 -88 -48 -86
rect -46 -88 -45 -86
rect -73 -95 -72 -93
rect -70 -95 -69 -93
rect -73 -96 -69 -95
rect -49 -94 -45 -88
rect -30 -84 -24 -83
rect -30 -86 -28 -84
rect -26 -86 -24 -84
rect -30 -90 -24 -86
rect -13 -84 0 -83
rect -13 -86 -6 -84
rect -4 -86 0 -84
rect -13 -87 0 -86
rect -47 -96 -45 -94
rect -31 -91 -17 -90
rect -31 -93 -30 -91
rect -28 -93 -17 -91
rect -31 -96 -17 -93
rect -13 -93 -9 -87
rect 11 -86 15 -75
rect 11 -88 12 -86
rect 14 -88 15 -86
rect -13 -95 -12 -93
rect -10 -95 -9 -93
rect -13 -96 -9 -95
rect -115 -102 -114 -100
rect -112 -102 -111 -100
rect -115 -104 -111 -102
rect -49 -104 -45 -96
rect 11 -94 15 -88
rect 13 -96 15 -94
rect 11 -104 15 -96
rect -135 -110 29 -109
rect -135 -112 -128 -110
rect -126 -112 -116 -110
rect -114 -112 -60 -110
rect -58 -112 -50 -110
rect -48 -112 0 -110
rect 2 -112 10 -110
rect 12 -112 29 -110
rect -135 -114 24 -112
rect 26 -114 29 -112
rect -135 -117 29 -114
rect -94 -123 -30 -122
rect -94 -125 -93 -123
rect -91 -125 -33 -123
rect -31 -125 -30 -123
rect -94 -126 -30 -125
rect 11 -126 15 -122
rect -131 -131 -19 -130
rect -131 -133 -130 -131
rect -128 -133 -85 -131
rect -83 -133 -22 -131
rect -20 -133 -19 -131
rect -131 -134 -19 -133
rect 11 -134 15 -130
rect -143 -139 -111 -138
rect -143 -141 -142 -139
rect -140 -141 -114 -139
rect -112 -141 -111 -139
rect -143 -142 -111 -141
rect -49 -139 -45 -138
rect -49 -141 -48 -139
rect -46 -141 -45 -139
rect -49 -142 -45 -141
rect 11 -139 15 -138
rect 11 -141 12 -139
rect 14 -141 15 -139
rect 11 -142 15 -141
rect -151 -147 -69 -146
rect -151 -149 -150 -147
rect -148 -149 -72 -147
rect -70 -149 -69 -147
rect -151 -150 -69 -149
rect -159 -155 -9 -154
rect -159 -157 -158 -155
rect -156 -157 -12 -155
rect -10 -157 -9 -155
rect -159 -158 -9 -157
<< alu2 >>
rect -49 67 -45 68
rect -49 65 -48 67
rect -46 65 -45 67
rect -143 59 -139 60
rect -143 57 -142 59
rect -140 57 -139 59
rect -159 51 -155 52
rect -159 49 -158 51
rect -156 49 -155 51
rect -159 -155 -155 49
rect -151 43 -147 44
rect -151 41 -150 43
rect -148 41 -147 43
rect -151 -147 -147 41
rect -143 -139 -139 57
rect -73 59 -69 60
rect -73 57 -72 59
rect -70 57 -69 59
rect -115 51 -111 52
rect -115 49 -114 51
rect -112 49 -111 51
rect -131 43 -127 44
rect -131 41 -130 43
rect -128 41 -127 43
rect -131 -4 -127 41
rect -115 12 -111 49
rect -85 51 -81 52
rect -85 49 -84 51
rect -82 49 -81 51
rect -115 10 -114 12
rect -112 10 -111 12
rect -115 8 -111 10
rect -94 35 -90 36
rect -94 33 -93 35
rect -91 33 -90 35
rect -131 -6 -130 -4
rect -128 -6 -127 -4
rect -131 -8 -127 -6
rect -94 -12 -90 33
rect -85 5 -81 49
rect -85 3 -84 5
rect -82 3 -81 5
rect -85 2 -81 3
rect -73 5 -69 57
rect -73 3 -72 5
rect -70 3 -69 5
rect -73 2 -69 3
rect -49 0 -45 65
rect 11 67 15 68
rect 11 65 12 67
rect 14 65 15 67
rect -13 59 -9 60
rect -13 57 -12 59
rect -10 57 -9 59
rect -23 43 -19 44
rect -23 41 -22 43
rect -20 41 -19 43
rect -34 35 -30 36
rect -34 33 -33 35
rect -31 33 -30 35
rect -34 19 -30 33
rect -49 -2 -48 0
rect -46 -2 -45 0
rect -49 -3 -45 -2
rect -35 4 -30 19
rect -35 3 -27 4
rect -35 1 -30 3
rect -28 1 -27 3
rect -35 0 -27 1
rect -94 -14 -93 -12
rect -91 -14 -90 -12
rect -94 -15 -90 -14
rect -83 -76 -79 -75
rect -83 -78 -82 -76
rect -80 -78 -79 -76
rect -131 -84 -127 -82
rect -131 -86 -130 -84
rect -128 -86 -127 -84
rect -131 -131 -127 -86
rect -95 -91 -87 -90
rect -95 -93 -90 -91
rect -88 -93 -87 -91
rect -95 -94 -87 -93
rect -131 -133 -130 -131
rect -128 -133 -127 -131
rect -131 -134 -127 -133
rect -115 -100 -111 -98
rect -115 -102 -114 -100
rect -112 -102 -111 -100
rect -143 -141 -142 -139
rect -140 -141 -139 -139
rect -143 -142 -139 -141
rect -115 -139 -111 -102
rect -95 -109 -90 -94
rect -83 -105 -79 -78
rect -49 -86 -45 -85
rect -49 -88 -48 -86
rect -46 -88 -45 -86
rect -94 -123 -90 -109
rect -94 -125 -93 -123
rect -91 -125 -90 -123
rect -94 -126 -90 -125
rect -86 -109 -79 -105
rect -73 -93 -69 -92
rect -73 -95 -72 -93
rect -70 -95 -69 -93
rect -86 -131 -82 -109
rect -86 -133 -85 -131
rect -83 -133 -82 -131
rect -86 -134 -82 -133
rect -115 -141 -114 -139
rect -112 -141 -111 -139
rect -115 -142 -111 -141
rect -151 -149 -150 -147
rect -148 -149 -147 -147
rect -151 -150 -147 -149
rect -73 -147 -69 -95
rect -49 -139 -45 -88
rect -35 -90 -30 0
rect -23 -12 -19 41
rect -13 5 -9 57
rect -13 3 -12 5
rect -10 3 -9 5
rect -13 2 -9 3
rect 11 0 15 65
rect 11 -2 12 0
rect 14 -2 15 0
rect 11 -3 15 -2
rect 22 24 29 27
rect 22 22 25 24
rect 27 22 29 24
rect -23 -14 -22 -12
rect -20 -14 -19 -12
rect -23 -15 -19 -14
rect -23 -76 -19 -75
rect -23 -78 -22 -76
rect -20 -78 -19 -76
rect -35 -91 -27 -90
rect -35 -93 -30 -91
rect -28 -93 -27 -91
rect -35 -94 -27 -93
rect -35 -122 -30 -94
rect -34 -123 -30 -122
rect -34 -125 -33 -123
rect -31 -125 -30 -123
rect -34 -126 -30 -125
rect -23 -131 -19 -78
rect 11 -86 15 -85
rect 11 -88 12 -86
rect 14 -88 15 -86
rect -23 -133 -22 -131
rect -20 -133 -19 -131
rect -23 -134 -19 -133
rect -13 -93 -9 -92
rect -13 -95 -12 -93
rect -10 -95 -9 -93
rect -49 -141 -48 -139
rect -46 -141 -45 -139
rect -49 -142 -45 -141
rect -73 -149 -72 -147
rect -70 -149 -69 -147
rect -73 -150 -69 -149
rect -159 -157 -158 -155
rect -156 -157 -155 -155
rect -159 -158 -155 -157
rect -13 -155 -9 -95
rect 11 -139 15 -88
rect 22 -112 29 22
rect 22 -114 24 -112
rect 26 -114 29 -112
rect 22 -117 29 -114
rect 11 -141 12 -139
rect 14 -141 15 -139
rect 11 -142 15 -141
rect -13 -157 -12 -155
rect -10 -157 -9 -155
rect -13 -158 -9 -157
<< ptie >>
rect -130 22 -112 24
rect -130 20 -128 22
rect -126 20 -116 22
rect -114 20 -112 22
rect -130 18 -112 20
rect -52 22 -46 24
rect -52 20 -50 22
rect -48 20 -46 22
rect -52 18 -46 20
rect 8 22 14 24
rect 8 20 10 22
rect 12 20 14 22
rect 8 18 14 20
rect -130 -110 -112 -108
rect -130 -112 -128 -110
rect -126 -112 -116 -110
rect -114 -112 -112 -110
rect -130 -114 -112 -112
rect -52 -110 -46 -108
rect -52 -112 -50 -110
rect -48 -112 -46 -110
rect -52 -114 -46 -112
rect 8 -110 14 -108
rect 8 -112 10 -110
rect 12 -112 14 -110
rect 8 -114 14 -112
<< ntie >>
rect -130 -38 -112 -36
rect -130 -40 -128 -38
rect -126 -40 -116 -38
rect -114 -40 -112 -38
rect -130 -42 -112 -40
rect -96 -38 -90 -36
rect -96 -40 -94 -38
rect -92 -40 -90 -38
rect -96 -42 -90 -40
rect -36 -38 -30 -36
rect -36 -40 -34 -38
rect -32 -40 -30 -38
rect -36 -42 -30 -40
rect -130 -50 -112 -48
rect -130 -52 -128 -50
rect -126 -52 -116 -50
rect -114 -52 -112 -50
rect -130 -54 -112 -52
rect -96 -50 -90 -48
rect -96 -52 -94 -50
rect -92 -52 -90 -50
rect -96 -54 -90 -52
rect -36 -50 -30 -48
rect -36 -52 -34 -50
rect -32 -52 -30 -50
rect -36 -54 -30 -52
<< nmos >>
rect -120 1 -118 10
rect -81 2 -79 15
rect -74 2 -72 15
rect -67 2 -65 15
rect -54 2 -52 11
rect -21 2 -19 15
rect -14 2 -12 15
rect -7 2 -5 15
rect 6 2 8 11
rect -120 -100 -118 -91
rect -81 -105 -79 -92
rect -74 -105 -72 -92
rect -67 -105 -65 -92
rect -54 -101 -52 -92
rect -21 -105 -19 -92
rect -14 -105 -12 -92
rect -7 -105 -5 -92
rect 6 -101 8 -92
<< pmos >>
rect -120 -29 -118 -11
rect -86 -30 -84 -17
rect -74 -31 -72 -18
rect -64 -31 -62 -18
rect -54 -31 -52 -13
rect -26 -30 -24 -17
rect -14 -31 -12 -18
rect -4 -31 -2 -18
rect 6 -31 8 -13
rect -120 -79 -118 -61
rect -86 -73 -84 -60
rect -74 -72 -72 -59
rect -64 -72 -62 -59
rect -54 -77 -52 -59
rect -26 -73 -24 -60
rect -14 -72 -12 -59
rect -4 -72 -2 -59
rect 6 -77 8 -59
<< polyct0 >>
rect -56 -6 -54 -4
rect 4 -6 6 -4
rect -56 -86 -54 -84
rect 4 -86 6 -84
<< polyct1 >>
rect -122 -6 -120 -4
rect -88 -6 -86 -4
rect -66 -6 -64 -4
rect -28 -6 -26 -4
rect -76 -13 -74 -11
rect -6 -6 -4 -4
rect -16 -13 -14 -11
rect -76 -79 -74 -77
rect -122 -86 -120 -84
rect -88 -86 -86 -84
rect -16 -79 -14 -77
rect -66 -86 -64 -84
rect -28 -86 -26 -84
rect -6 -86 -4 -84
<< ndifct0 >>
rect -86 11 -84 13
rect -129 6 -127 8
rect -26 11 -24 13
rect -129 -98 -127 -96
rect -86 -103 -84 -101
rect -26 -103 -24 -101
<< ndifct1 >>
rect -60 20 -58 22
rect 0 20 2 22
rect -115 3 -113 5
rect -49 4 -47 6
rect 11 4 13 6
rect -115 -95 -113 -93
rect -49 -96 -47 -94
rect 11 -96 13 -94
rect -60 -112 -58 -110
rect 0 -112 2 -110
<< ntiect1 >>
rect -128 -40 -126 -38
rect -116 -40 -114 -38
rect -94 -40 -92 -38
rect -34 -40 -32 -38
rect -128 -52 -126 -50
rect -116 -52 -114 -50
rect -94 -52 -92 -50
rect -34 -52 -32 -50
<< ptiect1 >>
rect -128 20 -126 22
rect -116 20 -114 22
rect -50 20 -48 22
rect 10 20 12 22
rect -128 -112 -126 -110
rect -116 -112 -114 -110
rect -50 -112 -48 -110
rect 10 -112 12 -110
<< pdifct0 >>
rect -126 -30 -124 -28
rect -91 -21 -89 -19
rect -91 -28 -89 -26
rect -69 -22 -67 -20
rect -69 -29 -67 -27
rect -59 -29 -57 -27
rect -31 -21 -29 -19
rect -31 -28 -29 -26
rect -9 -22 -7 -20
rect -9 -29 -7 -27
rect 1 -29 3 -27
rect -126 -62 -124 -60
rect -91 -64 -89 -62
rect -91 -71 -89 -69
rect -69 -63 -67 -61
rect -69 -70 -67 -68
rect -59 -63 -57 -61
rect -31 -64 -29 -62
rect -31 -71 -29 -69
rect -9 -63 -7 -61
rect -9 -70 -7 -68
rect 1 -63 3 -61
<< pdifct1 >>
rect -115 -15 -113 -13
rect -115 -22 -113 -20
rect -49 -17 -47 -15
rect -49 -24 -47 -22
rect 11 -17 13 -15
rect 11 -24 13 -22
rect -80 -40 -78 -38
rect -20 -40 -18 -38
rect -80 -52 -78 -50
rect -20 -52 -18 -50
rect -115 -70 -113 -68
rect -115 -77 -113 -75
rect -49 -68 -47 -66
rect -49 -75 -47 -73
rect 11 -68 13 -66
rect 11 -75 13 -73
<< alu0 >>
rect -130 8 -126 19
rect -130 6 -129 8
rect -127 6 -126 8
rect -88 13 -58 14
rect -88 11 -86 13
rect -84 11 -58 13
rect -88 10 -58 11
rect -130 4 -126 6
rect -116 1 -115 7
rect -62 6 -58 10
rect -116 -18 -115 -11
rect -62 2 -53 6
rect -50 2 -49 8
rect -28 13 2 14
rect -28 11 -26 13
rect -24 11 2 13
rect -28 10 2 11
rect -2 6 2 10
rect -57 -4 -53 2
rect -57 -6 -56 -4
rect -54 -6 -53 -4
rect -78 -11 -72 -10
rect -57 -11 -53 -6
rect -65 -15 -53 -11
rect -93 -19 -87 -18
rect -93 -21 -91 -19
rect -89 -21 -87 -19
rect -93 -26 -87 -21
rect -65 -18 -61 -15
rect -70 -20 -61 -18
rect -50 -19 -49 -13
rect -2 2 7 6
rect 10 2 11 8
rect 3 -4 7 2
rect 3 -6 4 -4
rect 6 -6 7 -4
rect -18 -11 -12 -10
rect 3 -11 7 -6
rect -5 -15 7 -11
rect -70 -22 -69 -20
rect -67 -22 -61 -20
rect -128 -28 -122 -27
rect -128 -30 -126 -28
rect -124 -30 -122 -28
rect -128 -37 -122 -30
rect -93 -28 -91 -26
rect -89 -27 -87 -26
rect -70 -27 -66 -22
rect -89 -28 -69 -27
rect -93 -29 -69 -28
rect -67 -29 -66 -27
rect -93 -31 -66 -29
rect -61 -27 -55 -26
rect -61 -29 -59 -27
rect -57 -29 -55 -27
rect -61 -37 -55 -29
rect -33 -19 -27 -18
rect -33 -21 -31 -19
rect -29 -21 -27 -19
rect -33 -26 -27 -21
rect -5 -18 -1 -15
rect -10 -20 -1 -18
rect 10 -19 11 -13
rect -10 -22 -9 -20
rect -7 -22 -1 -20
rect -33 -28 -31 -26
rect -29 -27 -27 -26
rect -10 -27 -6 -22
rect -29 -28 -9 -27
rect -33 -29 -9 -28
rect -7 -29 -6 -27
rect -33 -31 -6 -29
rect -1 -27 5 -26
rect -1 -29 1 -27
rect 3 -29 5 -27
rect -1 -37 5 -29
rect -128 -60 -122 -53
rect -128 -62 -126 -60
rect -124 -62 -122 -60
rect -128 -63 -122 -62
rect -93 -61 -66 -59
rect -93 -62 -69 -61
rect -93 -64 -91 -62
rect -89 -63 -69 -62
rect -67 -63 -66 -61
rect -89 -64 -87 -63
rect -93 -69 -87 -64
rect -93 -71 -91 -69
rect -89 -71 -87 -69
rect -93 -72 -87 -71
rect -116 -79 -115 -72
rect -70 -68 -66 -63
rect -61 -61 -55 -53
rect -61 -63 -59 -61
rect -57 -63 -55 -61
rect -61 -64 -55 -63
rect -70 -70 -69 -68
rect -67 -70 -61 -68
rect -70 -72 -61 -70
rect -65 -75 -61 -72
rect -130 -96 -126 -94
rect -130 -98 -129 -96
rect -127 -98 -126 -96
rect -116 -97 -115 -91
rect -65 -79 -53 -75
rect -50 -77 -49 -71
rect -33 -61 -6 -59
rect -33 -62 -9 -61
rect -33 -64 -31 -62
rect -29 -63 -9 -62
rect -7 -63 -6 -61
rect -29 -64 -27 -63
rect -33 -69 -27 -64
rect -33 -71 -31 -69
rect -29 -71 -27 -69
rect -33 -72 -27 -71
rect -10 -68 -6 -63
rect -1 -61 5 -53
rect -1 -63 1 -61
rect 3 -63 5 -61
rect -1 -64 5 -63
rect -10 -70 -9 -68
rect -7 -70 -1 -68
rect -10 -72 -1 -70
rect -5 -75 -1 -72
rect -78 -80 -72 -79
rect -57 -84 -53 -79
rect -57 -86 -56 -84
rect -54 -86 -53 -84
rect -130 -109 -126 -98
rect -57 -92 -53 -86
rect -5 -79 7 -75
rect 10 -77 11 -71
rect -18 -80 -12 -79
rect -62 -96 -53 -92
rect -62 -100 -58 -96
rect -50 -98 -49 -92
rect 3 -84 7 -79
rect 3 -86 4 -84
rect 6 -86 7 -84
rect 3 -92 7 -86
rect -2 -96 7 -92
rect -88 -101 -58 -100
rect -88 -103 -86 -101
rect -84 -103 -58 -101
rect -88 -104 -58 -103
rect -2 -100 2 -96
rect 10 -98 11 -92
rect -28 -101 2 -100
rect -28 -103 -26 -101
rect -24 -103 2 -101
rect -28 -104 2 -103
<< via1 >>
rect -48 65 -46 67
rect 12 65 14 67
rect -142 57 -140 59
rect -72 57 -70 59
rect -12 57 -10 59
rect -158 49 -156 51
rect -114 49 -112 51
rect -84 49 -82 51
rect -150 41 -148 43
rect -130 41 -128 43
rect -22 41 -20 43
rect -93 33 -91 35
rect -33 33 -31 35
rect 25 22 27 24
rect -114 10 -112 12
rect -130 -6 -128 -4
rect -84 3 -82 5
rect -72 3 -70 5
rect -93 -14 -91 -12
rect -30 1 -28 3
rect -12 3 -10 5
rect -48 -2 -46 0
rect -22 -14 -20 -12
rect 12 -2 14 0
rect -130 -86 -128 -84
rect -82 -78 -80 -76
rect -90 -93 -88 -91
rect -22 -78 -20 -76
rect -48 -88 -46 -86
rect -72 -95 -70 -93
rect -30 -93 -28 -91
rect 12 -88 14 -86
rect -12 -95 -10 -93
rect -114 -102 -112 -100
rect 24 -114 26 -112
rect -93 -125 -91 -123
rect -33 -125 -31 -123
rect -130 -133 -128 -131
rect -85 -133 -83 -131
rect -22 -133 -20 -131
rect -142 -141 -140 -139
rect -114 -141 -112 -139
rect -48 -141 -46 -139
rect 12 -141 14 -139
rect -150 -149 -148 -147
rect -72 -149 -70 -147
rect -158 -157 -156 -155
rect -12 -157 -10 -155
<< labels >>
rlabel alu1 -71 -49 -71 -49 4 vdd
rlabel alu1 -11 -49 -11 -49 4 vdd
rlabel alu1 -121 -49 -121 -49 4 vdd
rlabel via1 -92 -124 -92 -124 1 En
rlabel alu1 -71 -41 -71 -41 2 vdd
rlabel alu1 -11 -41 -11 -41 2 vdd
rlabel alu1 -121 -41 -121 -41 2 vdd
rlabel via1 -129 42 -129 42 1 A1
rlabel via1 -129 -132 -129 -132 1 A0
rlabel via1 13 66 13 66 5 Y2
rlabel via1 -47 66 -47 66 5 Y0
rlabel via1 -47 -140 -47 -140 1 Y3
rlabel via1 13 -140 13 -140 1 Y1
rlabel alu1 -104 23 -104 23 1 vss
rlabel alu1 -39 23 -39 23 1 vss
rlabel alu1 7 23 7 23 1 vss
rlabel alu1 -104 -113 -104 -113 1 vss
rlabel alu1 -54 -113 -54 -113 1 vss
rlabel alu1 6 -113 6 -113 1 vss
rlabel via1 -92 34 -92 34 1 En
<< end >>
