magic
tech scmos
timestamp 1607486678
<< ab >>
rect -179 -34 -157 38
rect -153 -34 -23 38
rect -21 -34 11 38
rect 14 -34 46 38
rect 49 -34 104 38
<< nwell >>
rect -184 -2 109 43
<< pwell >>
rect -184 -39 109 -2
<< poly >>
rect -168 22 -166 27
rect -142 22 -140 27
rect -120 23 -118 28
rect -10 32 -8 36
rect -3 32 -1 36
rect 25 32 27 36
rect 32 32 34 36
rect -108 24 -106 29
rect -98 24 -96 29
rect -88 24 -86 29
rect -168 1 -166 4
rect -142 1 -140 4
rect -120 1 -118 10
rect -108 8 -106 11
rect -112 6 -106 8
rect -112 4 -110 6
rect -108 4 -106 6
rect -112 2 -106 4
rect -172 -1 -166 1
rect -172 -3 -170 -1
rect -168 -3 -166 -1
rect -172 -5 -166 -3
rect -146 -1 -140 1
rect -146 -3 -144 -1
rect -142 -3 -140 -1
rect -146 -5 -140 -3
rect -124 -1 -118 1
rect -124 -3 -122 -1
rect -120 -3 -118 -1
rect -124 -5 -113 -3
rect -168 -8 -166 -5
rect -142 -8 -140 -5
rect -115 -9 -113 -5
rect -108 -9 -106 2
rect -98 1 -96 11
rect -66 23 -64 28
rect -54 24 -52 29
rect -44 24 -42 29
rect -34 24 -32 29
rect -88 1 -86 6
rect -66 1 -64 10
rect -54 8 -52 11
rect -58 6 -52 8
rect -58 4 -56 6
rect -54 4 -52 6
rect -58 2 -52 4
rect -102 -1 -96 1
rect -102 -3 -100 -1
rect -98 -3 -96 -1
rect -102 -5 -96 -3
rect -92 -1 -86 1
rect -92 -3 -90 -1
rect -88 -3 -86 -1
rect -92 -5 -86 -3
rect -70 -1 -64 1
rect -70 -3 -68 -1
rect -66 -3 -64 -1
rect -70 -5 -59 -3
rect -101 -9 -99 -5
rect -88 -9 -86 -5
rect -61 -9 -59 -5
rect -54 -9 -52 2
rect -44 1 -42 11
rect -34 1 -32 6
rect 60 23 62 28
rect 72 24 74 29
rect 82 24 84 29
rect 92 24 94 29
rect -48 -1 -42 1
rect -48 -3 -46 -1
rect -44 -3 -42 -1
rect -48 -5 -42 -3
rect -38 -1 -32 1
rect -38 -3 -36 -1
rect -34 -3 -32 -1
rect -10 -2 -8 4
rect -3 1 -1 4
rect -38 -5 -32 -3
rect -47 -9 -45 -5
rect -34 -9 -32 -5
rect -14 -4 -8 -2
rect -14 -6 -12 -4
rect -10 -6 -8 -4
rect -4 -1 2 1
rect -4 -3 -2 -1
rect 0 -3 2 -1
rect 25 -2 27 4
rect 32 1 34 4
rect 60 1 62 10
rect 72 8 74 11
rect 68 6 74 8
rect 68 4 70 6
rect 72 4 74 6
rect 68 2 74 4
rect -4 -5 2 -3
rect 21 -4 27 -2
rect -14 -8 -8 -6
rect -168 -22 -166 -17
rect -142 -22 -140 -17
rect -115 -27 -113 -22
rect -108 -27 -106 -22
rect -101 -27 -99 -22
rect -88 -23 -86 -18
rect -12 -11 -10 -8
rect -61 -27 -59 -22
rect -54 -27 -52 -22
rect -47 -27 -45 -22
rect -34 -23 -32 -18
rect -1 -14 1 -5
rect 21 -6 23 -4
rect 25 -6 27 -4
rect 31 -1 37 1
rect 31 -3 33 -1
rect 35 -3 37 -1
rect 31 -5 37 -3
rect 56 -1 62 1
rect 56 -3 58 -1
rect 60 -3 62 -1
rect 56 -5 67 -3
rect 21 -8 27 -6
rect 23 -11 25 -8
rect -12 -23 -10 -19
rect 34 -14 36 -5
rect 65 -9 67 -5
rect 72 -9 74 2
rect 82 1 84 11
rect 92 1 94 6
rect 78 -1 84 1
rect 78 -3 80 -1
rect 82 -3 84 -1
rect 78 -5 84 -3
rect 88 -1 94 1
rect 88 -3 90 -1
rect 92 -3 94 -1
rect 88 -5 94 -3
rect 79 -9 81 -5
rect 92 -9 94 -5
rect -1 -27 1 -22
rect 23 -23 25 -19
rect 34 -27 36 -22
rect 65 -27 67 -22
rect 72 -27 74 -22
rect 79 -27 81 -22
rect 92 -23 94 -18
<< ndif >>
rect -179 -13 -168 -8
rect -179 -15 -177 -13
rect -175 -15 -168 -13
rect -179 -17 -168 -15
rect -166 -10 -159 -8
rect -166 -12 -163 -10
rect -161 -12 -159 -10
rect -166 -14 -159 -12
rect -153 -13 -142 -8
rect -166 -17 -161 -14
rect -153 -15 -151 -13
rect -149 -15 -142 -13
rect -153 -17 -142 -15
rect -140 -10 -133 -8
rect -140 -12 -137 -10
rect -135 -12 -133 -10
rect -140 -14 -133 -12
rect -140 -17 -135 -14
rect -120 -16 -115 -9
rect -122 -18 -115 -16
rect -122 -20 -120 -18
rect -118 -20 -115 -18
rect -122 -22 -115 -20
rect -113 -22 -108 -9
rect -106 -22 -101 -9
rect -99 -18 -88 -9
rect -86 -11 -79 -9
rect -86 -13 -83 -11
rect -81 -13 -79 -11
rect -86 -15 -79 -13
rect -86 -18 -81 -15
rect -66 -16 -61 -9
rect -68 -18 -61 -16
rect -99 -22 -90 -18
rect -97 -27 -90 -22
rect -68 -20 -66 -18
rect -64 -20 -61 -18
rect -68 -22 -61 -20
rect -59 -22 -54 -9
rect -52 -22 -47 -9
rect -45 -18 -34 -9
rect -32 -11 -25 -9
rect -32 -13 -29 -11
rect -27 -13 -25 -11
rect -32 -15 -25 -13
rect -19 -15 -12 -11
rect -32 -18 -27 -15
rect -19 -17 -17 -15
rect -15 -17 -12 -15
rect -45 -22 -36 -18
rect -97 -29 -94 -27
rect -92 -29 -90 -27
rect -97 -31 -90 -29
rect -43 -27 -36 -22
rect -19 -19 -12 -17
rect -10 -14 -5 -11
rect -10 -18 -1 -14
rect -10 -19 -6 -18
rect -8 -20 -6 -19
rect -4 -20 -1 -18
rect -8 -22 -1 -20
rect 1 -22 9 -14
rect 16 -15 23 -11
rect 16 -17 18 -15
rect 20 -17 23 -15
rect 16 -19 23 -17
rect 25 -14 30 -11
rect 25 -18 34 -14
rect 25 -19 29 -18
rect -43 -29 -40 -27
rect -38 -29 -36 -27
rect -43 -31 -36 -29
rect 3 -27 9 -22
rect 27 -20 29 -19
rect 31 -20 34 -18
rect 27 -22 34 -20
rect 36 -22 44 -14
rect 60 -16 65 -9
rect 58 -18 65 -16
rect 58 -20 60 -18
rect 62 -20 65 -18
rect 58 -22 65 -20
rect 67 -22 72 -9
rect 74 -22 79 -9
rect 81 -18 92 -9
rect 94 -11 101 -9
rect 94 -13 97 -11
rect 99 -13 101 -11
rect 94 -15 101 -13
rect 94 -18 99 -15
rect 81 -22 90 -18
rect 3 -29 5 -27
rect 7 -29 9 -27
rect 3 -31 9 -29
rect 38 -27 44 -22
rect 83 -27 90 -22
rect 38 -29 40 -27
rect 42 -29 44 -27
rect 38 -31 44 -29
rect 83 -29 86 -27
rect 88 -29 90 -27
rect 83 -31 90 -29
<< pdif >>
rect -116 33 -110 35
rect -116 31 -114 33
rect -112 31 -110 33
rect -177 23 -170 25
rect -177 21 -174 23
rect -172 22 -170 23
rect -151 23 -144 25
rect -172 21 -168 22
rect -177 4 -168 21
rect -166 17 -161 22
rect -151 21 -148 23
rect -146 22 -144 23
rect -116 24 -110 31
rect -62 33 -56 35
rect -62 31 -60 33
rect -58 31 -56 33
rect -116 23 -108 24
rect -146 21 -142 22
rect -166 15 -159 17
rect -166 13 -163 15
rect -161 13 -159 15
rect -166 8 -159 13
rect -166 6 -163 8
rect -161 6 -159 8
rect -166 4 -159 6
rect -151 4 -142 21
rect -140 17 -135 22
rect -127 21 -120 23
rect -127 19 -125 21
rect -123 19 -120 21
rect -140 15 -133 17
rect -140 13 -137 15
rect -135 13 -133 15
rect -140 8 -133 13
rect -127 14 -120 19
rect -127 12 -125 14
rect -123 12 -120 14
rect -127 10 -120 12
rect -118 11 -108 23
rect -106 22 -98 24
rect -106 20 -103 22
rect -101 20 -98 22
rect -106 15 -98 20
rect -106 13 -103 15
rect -101 13 -98 15
rect -106 11 -98 13
rect -96 22 -88 24
rect -96 20 -93 22
rect -91 20 -88 22
rect -96 11 -88 20
rect -118 10 -113 11
rect -140 6 -137 8
rect -135 6 -133 8
rect -140 4 -133 6
rect -94 6 -88 11
rect -86 19 -81 24
rect -62 24 -56 31
rect -19 30 -10 32
rect -19 28 -17 30
rect -15 28 -10 30
rect -62 23 -54 24
rect -73 21 -66 23
rect -73 19 -71 21
rect -69 19 -66 21
rect -86 17 -79 19
rect -86 15 -83 17
rect -81 15 -79 17
rect -86 10 -79 15
rect -73 14 -66 19
rect -73 12 -71 14
rect -69 12 -66 14
rect -73 10 -66 12
rect -64 11 -54 23
rect -52 22 -44 24
rect -52 20 -49 22
rect -47 20 -44 22
rect -52 15 -44 20
rect -52 13 -49 15
rect -47 13 -44 15
rect -52 11 -44 13
rect -42 22 -34 24
rect -42 20 -39 22
rect -37 20 -34 22
rect -42 11 -34 20
rect -64 10 -59 11
rect -86 8 -83 10
rect -81 8 -79 10
rect -86 6 -79 8
rect -40 6 -34 11
rect -32 19 -27 24
rect -19 23 -10 28
rect -19 21 -17 23
rect -15 21 -10 23
rect -32 17 -25 19
rect -32 15 -29 17
rect -27 15 -25 17
rect -32 10 -25 15
rect -32 8 -29 10
rect -27 8 -25 10
rect -32 6 -25 8
rect -19 4 -10 21
rect -8 4 -3 32
rect -1 25 4 32
rect 16 30 25 32
rect 16 28 18 30
rect 20 28 25 30
rect -1 23 6 25
rect -1 21 2 23
rect 4 21 6 23
rect -1 16 6 21
rect -1 14 2 16
rect 4 14 6 16
rect -1 12 6 14
rect 16 23 25 28
rect 16 21 18 23
rect 20 21 25 23
rect -1 4 4 12
rect 16 4 25 21
rect 27 4 32 32
rect 34 25 39 32
rect 64 33 70 35
rect 64 31 66 33
rect 68 31 70 33
rect 34 23 41 25
rect 64 24 70 31
rect 64 23 72 24
rect 34 21 37 23
rect 39 21 41 23
rect 34 16 41 21
rect 34 14 37 16
rect 39 14 41 16
rect 34 12 41 14
rect 53 21 60 23
rect 53 19 55 21
rect 57 19 60 21
rect 53 14 60 19
rect 53 12 55 14
rect 57 12 60 14
rect 34 4 39 12
rect 53 10 60 12
rect 62 11 72 23
rect 74 22 82 24
rect 74 20 77 22
rect 79 20 82 22
rect 74 15 82 20
rect 74 13 77 15
rect 79 13 82 15
rect 74 11 82 13
rect 84 22 92 24
rect 84 20 87 22
rect 89 20 92 22
rect 84 11 92 20
rect 62 10 67 11
rect 86 6 92 11
rect 94 19 99 24
rect 94 17 101 19
rect 94 15 97 17
rect 99 15 101 17
rect 94 10 101 15
rect 94 8 97 10
rect 99 8 101 10
rect 94 6 101 8
<< alu1 >>
rect -179 33 106 38
rect -179 31 -176 33
rect -174 31 -164 33
rect -162 31 -150 33
rect -148 31 -138 33
rect -136 31 -128 33
rect -126 31 -114 33
rect -112 31 -74 33
rect -72 31 -60 33
rect -58 31 52 33
rect 54 31 66 33
rect 68 31 106 33
rect -179 30 106 31
rect -171 15 -159 17
rect -171 13 -163 15
rect -161 13 -159 15
rect -171 11 -159 13
rect -145 15 -133 17
rect -145 13 -137 15
rect -135 13 -133 15
rect -145 11 -133 13
rect -163 8 -159 11
rect -161 6 -159 8
rect -179 -1 -167 1
rect -179 -3 -177 -1
rect -175 -3 -170 -1
rect -168 -3 -167 -1
rect -179 -5 -167 -3
rect -171 -13 -167 -5
rect -163 -4 -159 6
rect -137 8 -133 11
rect -116 8 -110 16
rect -84 17 -79 25
rect -84 16 -83 17
rect -92 15 -83 16
rect -81 15 -79 17
rect -92 12 -79 15
rect -135 6 -133 8
rect -163 -6 -162 -4
rect -160 -6 -159 -4
rect -153 -1 -141 1
rect -153 -3 -152 -1
rect -150 -3 -144 -1
rect -142 -3 -141 -1
rect -153 -5 -141 -3
rect -163 -10 -159 -6
rect -161 -12 -159 -10
rect -163 -21 -159 -12
rect -145 -13 -141 -5
rect -137 -4 -133 6
rect -124 7 -102 8
rect -124 5 -115 7
rect -113 6 -102 7
rect -113 5 -110 6
rect -124 4 -110 5
rect -108 4 -102 6
rect -83 10 -79 12
rect -81 8 -79 10
rect -62 8 -56 16
rect -30 17 -25 25
rect 0 23 6 24
rect 0 21 2 23
rect 4 21 6 23
rect -30 16 -29 17
rect -38 15 -29 16
rect -27 15 -25 17
rect -38 12 -25 15
rect 0 17 6 21
rect 35 23 41 24
rect 35 21 37 23
rect 39 21 41 23
rect 35 17 41 21
rect 0 16 9 17
rect 0 14 2 16
rect 4 14 9 16
rect 0 13 9 14
rect 35 16 44 17
rect 35 14 37 16
rect 39 14 44 16
rect 35 13 44 14
rect -137 -6 -136 -4
rect -134 -6 -133 -4
rect -137 -10 -133 -6
rect -135 -12 -133 -10
rect -137 -21 -133 -12
rect -124 -1 -118 0
rect -124 -3 -122 -1
rect -120 -3 -118 -1
rect -124 -7 -118 -3
rect -107 -1 -94 0
rect -107 -3 -100 -1
rect -98 -3 -94 -1
rect -107 -4 -94 -3
rect -124 -10 -111 -7
rect -124 -12 -123 -10
rect -121 -12 -111 -10
rect -124 -13 -111 -12
rect -107 -8 -103 -4
rect -107 -10 -106 -8
rect -104 -10 -103 -8
rect -83 -3 -79 8
rect -70 7 -48 8
rect -70 5 -61 7
rect -59 6 -48 7
rect -59 5 -56 6
rect -70 4 -56 5
rect -54 4 -48 6
rect -29 10 -25 12
rect -27 8 -25 10
rect -83 -5 -82 -3
rect -80 -5 -79 -3
rect -107 -13 -103 -10
rect -83 -11 -79 -5
rect -81 -13 -79 -11
rect -70 -1 -64 0
rect -70 -3 -68 -1
rect -66 -3 -64 -1
rect -70 -7 -64 -3
rect -53 -1 -40 0
rect -53 -3 -46 -1
rect -44 -3 -40 -1
rect -53 -4 -40 -3
rect -70 -10 -57 -7
rect -70 -12 -69 -10
rect -67 -12 -57 -10
rect -70 -13 -57 -12
rect -53 -8 -49 -4
rect -53 -10 -52 -8
rect -50 -10 -49 -8
rect -29 -3 -25 8
rect -11 5 -7 9
rect -11 4 1 5
rect -11 2 -2 4
rect 0 2 1 4
rect -11 1 1 2
rect -29 -5 -28 -3
rect -26 -5 -25 -3
rect -53 -13 -49 -10
rect -83 -21 -79 -13
rect -29 -11 -25 -5
rect -19 -3 -15 1
rect -3 -1 1 1
rect -3 -3 -2 -1
rect 0 -3 1 -1
rect -19 -4 -7 -3
rect -19 -6 -18 -4
rect -16 -6 -12 -4
rect -10 -6 -7 -4
rect -3 -5 1 -3
rect -19 -7 -7 -6
rect -27 -13 -25 -11
rect -11 -13 -7 -7
rect 5 -9 9 13
rect 24 5 28 9
rect 24 4 36 5
rect 24 2 29 4
rect 31 2 36 4
rect 24 1 36 2
rect 16 -3 20 1
rect 32 -1 36 1
rect 32 -3 33 -1
rect 35 -3 36 -1
rect 16 -4 28 -3
rect 16 -6 17 -4
rect 19 -6 23 -4
rect 25 -6 28 -4
rect 32 -5 36 -3
rect 16 -7 28 -6
rect 5 -11 6 -9
rect 8 -11 9 -9
rect -29 -21 -25 -13
rect 5 -15 9 -11
rect 24 -13 28 -7
rect 40 -11 44 13
rect 64 8 70 16
rect 96 17 101 25
rect 96 16 97 17
rect 88 15 97 16
rect 99 15 101 17
rect 88 12 101 15
rect 56 7 78 8
rect 56 5 65 7
rect 67 6 78 7
rect 67 5 70 6
rect 56 4 70 5
rect 72 4 78 6
rect 97 10 101 12
rect 99 8 101 10
rect 40 -13 41 -11
rect 43 -13 44 -11
rect 56 -1 62 0
rect 56 -3 58 -1
rect 60 -3 62 -1
rect 56 -7 62 -3
rect 73 -1 86 0
rect 73 -3 80 -1
rect 82 -3 86 -1
rect 73 -4 86 -3
rect 56 -10 69 -7
rect 56 -12 57 -10
rect 59 -12 69 -10
rect 56 -13 69 -12
rect 73 -9 77 -4
rect 97 -7 101 8
rect 97 -9 98 -7
rect 100 -9 101 -7
rect 73 -11 74 -9
rect 76 -11 77 -9
rect 73 -13 77 -11
rect -3 -17 9 -15
rect -8 -18 9 -17
rect -8 -20 -6 -18
rect -4 -20 9 -18
rect -8 -21 9 -20
rect 40 -15 44 -13
rect 32 -17 44 -15
rect 97 -11 101 -9
rect 99 -13 101 -11
rect 27 -18 44 -17
rect 27 -20 29 -18
rect 31 -20 44 -18
rect 27 -21 44 -20
rect 97 -21 101 -13
rect -179 -27 106 -26
rect -179 -29 -176 -27
rect -174 -29 -164 -27
rect -162 -29 -150 -27
rect -148 -29 -138 -27
rect -136 -29 -94 -27
rect -92 -29 -84 -27
rect -82 -29 -40 -27
rect -38 -29 -30 -27
rect -28 -29 -16 -27
rect -14 -29 5 -27
rect 7 -29 19 -27
rect 21 -29 40 -27
rect 42 -29 86 -27
rect 88 -29 96 -27
rect 98 -29 106 -27
rect -179 -34 106 -29
rect -163 -40 -120 -39
rect -163 -42 -162 -40
rect -160 -42 -123 -40
rect -121 -42 -120 -40
rect -163 -43 -120 -42
rect -29 -40 -15 -39
rect -29 -42 -28 -40
rect -26 -42 -18 -40
rect -16 -42 -15 -40
rect -29 -43 -15 -42
rect 5 -40 20 -39
rect 5 -42 6 -40
rect 8 -42 17 -40
rect 19 -42 20 -40
rect 5 -43 20 -42
rect 28 -40 32 -39
rect 28 -42 29 -40
rect 31 -42 32 -40
rect 28 -43 32 -42
rect -178 -48 -66 -47
rect -178 -50 -177 -48
rect -175 -50 -69 -48
rect -67 -50 -66 -48
rect -178 -51 -66 -50
rect -3 -48 60 -47
rect -3 -50 -2 -48
rect 0 -50 41 -48
rect 43 -50 57 -48
rect 59 -50 60 -48
rect -3 -51 60 -50
rect -137 -56 -58 -55
rect -137 -58 -136 -56
rect -134 -58 -115 -56
rect -113 -58 -61 -56
rect -59 -58 -58 -56
rect -137 -59 -58 -58
rect -83 -64 32 -63
rect -83 -66 -82 -64
rect -80 -66 29 -64
rect 31 -66 32 -64
rect -83 -67 32 -66
rect -153 -72 68 -71
rect -153 -74 -152 -72
rect -150 -74 65 -72
rect 67 -74 68 -72
rect -153 -75 68 -74
rect -107 -80 77 -79
rect -107 -82 -106 -80
rect -104 -82 -52 -80
rect -50 -82 74 -80
rect 76 -82 77 -80
rect -107 -83 77 -82
<< alu2 >>
rect -116 7 -112 8
rect -116 5 -115 7
rect -113 5 -112 7
rect -178 -1 -174 0
rect -178 -3 -177 -1
rect -175 -3 -174 -1
rect -153 -1 -149 1
rect -153 -3 -152 -1
rect -150 -3 -149 -1
rect -178 -48 -174 -3
rect -163 -4 -159 -3
rect -163 -6 -162 -4
rect -160 -6 -159 -4
rect -163 -40 -159 -6
rect -163 -42 -162 -40
rect -160 -42 -159 -40
rect -163 -43 -159 -42
rect -178 -50 -177 -48
rect -175 -50 -174 -48
rect -178 -51 -174 -50
rect -153 -72 -149 -3
rect -137 -4 -133 -3
rect -137 -6 -136 -4
rect -134 -6 -133 -4
rect -137 -56 -133 -6
rect -124 -10 -120 -9
rect -124 -12 -123 -10
rect -121 -12 -120 -10
rect -124 -40 -120 -12
rect -124 -42 -123 -40
rect -121 -42 -120 -40
rect -124 -43 -120 -42
rect -137 -58 -136 -56
rect -134 -58 -133 -56
rect -137 -59 -133 -58
rect -116 -56 -112 5
rect -62 7 -58 8
rect -62 5 -61 7
rect -59 5 -58 7
rect 64 7 68 8
rect 64 5 65 7
rect 67 5 68 7
rect -83 -3 -79 -2
rect -83 -5 -82 -3
rect -80 -5 -79 -3
rect -116 -58 -115 -56
rect -113 -58 -112 -56
rect -116 -59 -112 -58
rect -107 -8 -103 -7
rect -107 -10 -106 -8
rect -104 -10 -103 -8
rect -153 -74 -152 -72
rect -150 -74 -149 -72
rect -153 -75 -149 -74
rect -107 -80 -103 -10
rect -83 -64 -79 -5
rect -70 -10 -66 -9
rect -70 -12 -69 -10
rect -67 -12 -66 -10
rect -70 -48 -66 -12
rect -70 -50 -69 -48
rect -67 -50 -66 -48
rect -70 -51 -66 -50
rect -62 -56 -58 5
rect -3 4 1 5
rect -3 2 -2 4
rect 0 2 1 4
rect -29 -3 -25 -2
rect -29 -5 -28 -3
rect -26 -5 -25 -3
rect -62 -58 -61 -56
rect -59 -58 -58 -56
rect -62 -59 -58 -58
rect -53 -8 -49 -7
rect -53 -10 -52 -8
rect -50 -10 -49 -8
rect -83 -66 -82 -64
rect -80 -66 -79 -64
rect -83 -67 -79 -66
rect -107 -82 -106 -80
rect -104 -82 -103 -80
rect -107 -83 -103 -82
rect -53 -80 -49 -10
rect -29 -40 -25 -5
rect -29 -42 -28 -40
rect -26 -42 -25 -40
rect -29 -43 -25 -42
rect -19 -4 -15 -3
rect -19 -6 -18 -4
rect -16 -6 -15 -4
rect -19 -40 -15 -6
rect -19 -42 -18 -40
rect -16 -42 -15 -40
rect -19 -43 -15 -42
rect -3 -48 1 2
rect 28 4 32 5
rect 28 2 29 4
rect 31 2 32 4
rect 16 -4 20 -3
rect 16 -6 17 -4
rect 19 -6 20 -4
rect 5 -9 9 -8
rect 5 -11 6 -9
rect 8 -11 9 -9
rect 5 -40 9 -11
rect 5 -42 6 -40
rect 8 -42 9 -40
rect 5 -43 9 -42
rect 16 -40 20 -6
rect 16 -42 17 -40
rect 19 -42 20 -40
rect 16 -43 20 -42
rect 28 -40 32 2
rect 56 -10 60 -9
rect 28 -42 29 -40
rect 31 -42 32 -40
rect -3 -50 -2 -48
rect 0 -50 1 -48
rect -3 -51 1 -50
rect 28 -64 32 -42
rect 40 -11 44 -10
rect 40 -13 41 -11
rect 43 -13 44 -11
rect 40 -48 44 -13
rect 40 -50 41 -48
rect 43 -50 44 -48
rect 40 -51 44 -50
rect 56 -12 57 -10
rect 59 -12 60 -10
rect 56 -48 60 -12
rect 56 -50 57 -48
rect 59 -50 60 -48
rect 56 -51 60 -50
rect 28 -66 29 -64
rect 31 -66 32 -64
rect 28 -67 32 -66
rect 64 -72 68 5
rect 64 -74 65 -72
rect 67 -74 68 -72
rect 64 -75 68 -74
rect 73 -9 77 -7
rect 73 -11 74 -9
rect 76 -11 77 -9
rect -53 -82 -52 -80
rect -50 -82 -49 -80
rect -53 -83 -49 -82
rect 73 -80 77 -11
rect 83 -34 87 0
rect 97 -7 101 -6
rect 97 -9 98 -7
rect 100 -9 101 -7
rect 97 -53 101 -9
rect 73 -82 74 -80
rect 76 -82 77 -80
rect 73 -83 77 -82
<< ptie >>
rect -178 -27 -160 -25
rect -178 -29 -176 -27
rect -174 -29 -164 -27
rect -162 -29 -160 -27
rect -178 -31 -160 -29
rect -152 -27 -134 -25
rect -152 -29 -150 -27
rect -148 -29 -138 -27
rect -136 -29 -134 -27
rect -152 -31 -134 -29
rect -86 -27 -80 -25
rect -86 -29 -84 -27
rect -82 -29 -80 -27
rect -86 -31 -80 -29
rect -32 -27 -26 -25
rect -32 -29 -30 -27
rect -28 -29 -26 -27
rect -32 -31 -26 -29
rect -18 -27 -12 -25
rect -18 -29 -16 -27
rect -14 -29 -12 -27
rect -18 -31 -12 -29
rect 17 -27 23 -25
rect 17 -29 19 -27
rect 21 -29 23 -27
rect 17 -31 23 -29
rect 94 -27 100 -25
rect 94 -29 96 -27
rect 98 -29 100 -27
rect 94 -31 100 -29
<< ntie >>
rect -178 33 -160 35
rect -178 31 -176 33
rect -174 31 -164 33
rect -162 31 -160 33
rect -178 29 -160 31
rect -152 33 -134 35
rect -152 31 -150 33
rect -148 31 -138 33
rect -136 31 -134 33
rect -152 29 -134 31
rect -130 33 -124 35
rect -130 31 -128 33
rect -126 31 -124 33
rect -130 29 -124 31
rect -76 33 -70 35
rect -76 31 -74 33
rect -72 31 -70 33
rect -76 29 -70 31
rect 50 33 56 35
rect 50 31 52 33
rect 54 31 56 33
rect 50 29 56 31
<< nmos >>
rect -168 -17 -166 -8
rect -142 -17 -140 -8
rect -115 -22 -113 -9
rect -108 -22 -106 -9
rect -101 -22 -99 -9
rect -88 -18 -86 -9
rect -61 -22 -59 -9
rect -54 -22 -52 -9
rect -47 -22 -45 -9
rect -34 -18 -32 -9
rect -12 -19 -10 -11
rect -1 -22 1 -14
rect 23 -19 25 -11
rect 34 -22 36 -14
rect 65 -22 67 -9
rect 72 -22 74 -9
rect 79 -22 81 -9
rect 92 -18 94 -9
<< pmos >>
rect -168 4 -166 22
rect -142 4 -140 22
rect -120 10 -118 23
rect -108 11 -106 24
rect -98 11 -96 24
rect -88 6 -86 24
rect -66 10 -64 23
rect -54 11 -52 24
rect -44 11 -42 24
rect -34 6 -32 24
rect -10 4 -8 32
rect -3 4 -1 32
rect 25 4 27 32
rect 32 4 34 32
rect 60 10 62 23
rect 72 11 74 24
rect 82 11 84 24
rect 92 6 94 24
<< polyct0 >>
rect -90 -3 -88 -1
rect -36 -3 -34 -1
rect 90 -3 92 -1
<< polyct1 >>
rect -110 4 -108 6
rect -170 -3 -168 -1
rect -144 -3 -142 -1
rect -122 -3 -120 -1
rect -56 4 -54 6
rect -100 -3 -98 -1
rect -68 -3 -66 -1
rect -46 -3 -44 -1
rect -12 -6 -10 -4
rect -2 -3 0 -1
rect 70 4 72 6
rect 23 -6 25 -4
rect 33 -3 35 -1
rect 58 -3 60 -1
rect 80 -3 82 -1
<< ndifct0 >>
rect -177 -15 -175 -13
rect -151 -15 -149 -13
rect -120 -20 -118 -18
rect -66 -20 -64 -18
rect -17 -17 -15 -15
rect 18 -17 20 -15
rect 60 -20 62 -18
<< ndifct1 >>
rect -163 -12 -161 -10
rect -137 -12 -135 -10
rect -83 -13 -81 -11
rect -29 -13 -27 -11
rect -94 -29 -92 -27
rect -6 -20 -4 -18
rect -40 -29 -38 -27
rect 29 -20 31 -18
rect 97 -13 99 -11
rect 5 -29 7 -27
rect 40 -29 42 -27
rect 86 -29 88 -27
<< ntiect1 >>
rect -176 31 -174 33
rect -164 31 -162 33
rect -150 31 -148 33
rect -138 31 -136 33
rect -128 31 -126 33
rect -74 31 -72 33
rect 52 31 54 33
<< ptiect1 >>
rect -176 -29 -174 -27
rect -164 -29 -162 -27
rect -150 -29 -148 -27
rect -138 -29 -136 -27
rect -84 -29 -82 -27
rect -30 -29 -28 -27
rect -16 -29 -14 -27
rect 19 -29 21 -27
rect 96 -29 98 -27
<< pdifct0 >>
rect -174 21 -172 23
rect -148 21 -146 23
rect -125 19 -123 21
rect -125 12 -123 14
rect -103 20 -101 22
rect -103 13 -101 15
rect -93 20 -91 22
rect -17 28 -15 30
rect -71 19 -69 21
rect -71 12 -69 14
rect -49 20 -47 22
rect -49 13 -47 15
rect -39 20 -37 22
rect -17 21 -15 23
rect 18 28 20 30
rect 18 21 20 23
rect 55 19 57 21
rect 55 12 57 14
rect 77 20 79 22
rect 77 13 79 15
rect 87 20 89 22
<< pdifct1 >>
rect -114 31 -112 33
rect -60 31 -58 33
rect -163 13 -161 15
rect -163 6 -161 8
rect -137 13 -135 15
rect -137 6 -135 8
rect -83 15 -81 17
rect -83 8 -81 10
rect -29 15 -27 17
rect -29 8 -27 10
rect 2 21 4 23
rect 2 14 4 16
rect 66 31 68 33
rect 37 21 39 23
rect 37 14 39 16
rect 97 15 99 17
rect 97 8 99 10
<< alu0 >>
rect -176 23 -170 30
rect -176 21 -174 23
rect -172 21 -170 23
rect -176 20 -170 21
rect -150 23 -144 30
rect -150 21 -148 23
rect -146 21 -144 23
rect -150 20 -144 21
rect -127 22 -100 24
rect -127 21 -103 22
rect -127 19 -125 21
rect -123 20 -103 21
rect -101 20 -100 22
rect -123 19 -121 20
rect -127 14 -121 19
rect -127 12 -125 14
rect -123 12 -121 14
rect -127 11 -121 12
rect -164 4 -163 11
rect -178 -13 -174 -11
rect -138 4 -137 11
rect -104 15 -100 20
rect -95 22 -89 30
rect -95 20 -93 22
rect -91 20 -89 22
rect -95 19 -89 20
rect -104 13 -103 15
rect -101 13 -95 15
rect -104 11 -95 13
rect -99 8 -95 11
rect -178 -15 -177 -13
rect -175 -15 -174 -13
rect -164 -14 -163 -8
rect -178 -26 -174 -15
rect -152 -13 -148 -11
rect -99 4 -87 8
rect -84 6 -83 12
rect -73 22 -46 24
rect -73 21 -49 22
rect -73 19 -71 21
rect -69 20 -49 21
rect -47 20 -46 22
rect -69 19 -67 20
rect -73 14 -67 19
rect -73 12 -71 14
rect -69 12 -67 14
rect -73 11 -67 12
rect -50 15 -46 20
rect -41 22 -35 30
rect -18 28 -17 30
rect -15 28 -14 30
rect -41 20 -39 22
rect -37 20 -35 22
rect -41 19 -35 20
rect -18 23 -14 28
rect 17 28 18 30
rect 20 28 21 30
rect -18 21 -17 23
rect -15 21 -14 23
rect -18 19 -14 21
rect -50 13 -49 15
rect -47 13 -41 15
rect -50 11 -41 13
rect 17 23 21 28
rect 17 21 18 23
rect 20 21 21 23
rect 17 19 21 21
rect 53 22 80 24
rect 53 21 77 22
rect 53 19 55 21
rect 57 20 77 21
rect 79 20 80 22
rect 57 19 59 20
rect -45 8 -41 11
rect -112 3 -106 4
rect -152 -15 -151 -13
rect -149 -15 -148 -13
rect -138 -14 -137 -8
rect -152 -26 -148 -15
rect -91 -1 -87 4
rect -91 -3 -90 -1
rect -88 -3 -87 -1
rect -91 -9 -87 -3
rect -45 4 -33 8
rect -30 6 -29 12
rect -58 3 -52 4
rect -96 -13 -87 -9
rect -96 -17 -92 -13
rect -84 -15 -83 -9
rect -37 -1 -33 4
rect -37 -3 -36 -1
rect -34 -3 -33 -1
rect -37 -9 -33 -3
rect -42 -13 -33 -9
rect -122 -18 -92 -17
rect -122 -20 -120 -18
rect -118 -20 -92 -18
rect -122 -21 -92 -20
rect -42 -17 -38 -13
rect -30 -15 -29 -9
rect -68 -18 -38 -17
rect -68 -20 -66 -18
rect -64 -20 -38 -18
rect -68 -21 -38 -20
rect -18 -15 -14 -13
rect 53 14 59 19
rect 53 12 55 14
rect 57 12 59 14
rect 53 11 59 12
rect 76 15 80 20
rect 85 22 91 30
rect 85 20 87 22
rect 89 20 91 22
rect 85 19 91 20
rect 76 13 77 15
rect 79 13 85 15
rect 76 11 85 13
rect 81 8 85 11
rect 81 4 93 8
rect 96 6 97 12
rect 68 3 74 4
rect 89 -1 93 4
rect 89 -3 90 -1
rect 92 -3 93 -1
rect 89 -9 93 -3
rect 84 -13 93 -9
rect -18 -17 -17 -15
rect -15 -17 -14 -15
rect -18 -26 -14 -17
rect 17 -15 21 -13
rect 17 -17 18 -15
rect 20 -17 21 -15
rect 84 -17 88 -13
rect 96 -15 97 -9
rect 17 -26 21 -17
rect 58 -18 88 -17
rect 58 -20 60 -18
rect 62 -20 88 -18
rect 58 -21 88 -20
<< via1 >>
rect -177 -3 -175 -1
rect -162 -6 -160 -4
rect -152 -3 -150 -1
rect -115 5 -113 7
rect -136 -6 -134 -4
rect -123 -12 -121 -10
rect -106 -10 -104 -8
rect -61 5 -59 7
rect -82 -5 -80 -3
rect -69 -12 -67 -10
rect -52 -10 -50 -8
rect -2 2 0 4
rect -28 -5 -26 -3
rect -18 -6 -16 -4
rect 29 2 31 4
rect 17 -6 19 -4
rect 6 -11 8 -9
rect 65 5 67 7
rect 41 -13 43 -11
rect 57 -12 59 -10
rect 98 -9 100 -7
rect 74 -11 76 -9
rect -162 -42 -160 -40
rect -123 -42 -121 -40
rect -28 -42 -26 -40
rect -18 -42 -16 -40
rect 6 -42 8 -40
rect 17 -42 19 -40
rect 29 -42 31 -40
rect -177 -50 -175 -48
rect -69 -50 -67 -48
rect -2 -50 0 -48
rect 41 -50 43 -48
rect 57 -50 59 -48
rect -136 -58 -134 -56
rect -115 -58 -113 -56
rect -61 -58 -59 -56
rect -82 -66 -80 -64
rect 29 -66 31 -64
rect -152 -74 -150 -72
rect 65 -74 67 -72
rect -106 -82 -104 -80
rect -52 -82 -50 -80
rect 74 -82 76 -80
<< labels >>
rlabel alu1 75 -30 75 -30 4 vss
rlabel alu1 75 34 75 34 4 vdd
rlabel alu1 -51 -30 -51 -30 4 vss
rlabel alu1 -51 34 -51 34 4 vdd
rlabel alu1 -105 34 -105 34 4 vdd
rlabel alu1 -105 -30 -105 -30 4 vss
rlabel alu1 -169 34 -169 34 4 vdd
rlabel alu1 -169 -30 -169 -30 4 vss
rlabel alu1 -143 -30 -143 -30 4 vss
rlabel alu1 -143 34 -143 34 4 vdd
rlabel via1 -176 -49 -176 -49 1 Input
rlabel alu2 99 -49 99 -49 1 Output
rlabel via1 -151 -73 -151 -73 1 RorW
rlabel via1 -105 -81 -105 -81 1 Select
rlabel via1 30 -41 30 -41 1 R
rlabel via1 -17 -41 -17 -41 1 S
rlabel via1 42 -49 42 -49 1 Q
rlabel via1 7 -41 7 -41 1 Q_bar
rlabel alu1 30 -30 30 -30 4 vss
rlabel alu1 30 34 30 34 4 vdd
rlabel alu1 -5 34 -5 34 4 vdd
rlabel alu1 -5 -30 -5 -30 4 vss
<< end >>
